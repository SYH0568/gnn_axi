`timescale 1 ns / 1 ps

module AESL_deadlock_report_unit #( parameter PROC_NUM = 4 ) (
    input reset,
    input clock,
    input [PROC_NUM - 1:0] dl_in_vec,
    output dl_detect_out,
    output reg [PROC_NUM - 1:0] origin,
    output token_clear);
   
    // FSM states
    localparam ST_IDLE = 2'b0;
    localparam ST_DL_DETECTED = 2'b1;
    localparam ST_DL_REPORT = 2'b10;

    reg [1:0] CS_fsm;
    reg [1:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg) begin
        NS_fsm = CS_fsm;
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = |dl_detect_reg;

    // dl_done_reg record the cycles has been reported
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    always @ (CS_fsm or dl_detect_reg or dl_done_reg) begin
        origin = 'b0;
        if (CS_fsm == ST_DL_DETECTED) begin
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_detect_reg[i] & ~dl_done_reg[i] & ~(|origin)) begin
                    origin = 'b1 << i;
                end
            end
        end
    end
    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [344:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "example.Block_proc_U0";
                end
                1 : begin
                    proc_path = "example.clone_vector_3_U0";
                end
                2 : begin
                    proc_path = "example.clone_vector_1_U0";
                end
                3 : begin
                    proc_path = "example.clone_vector_U0";
                end
                4 : begin
                    proc_path = "example.Loop_edge_choose_ver_1_U0";
                end
                5 : begin
                    proc_path = "example.Loop_edge_compute_lo_1_U0";
                end
                6 : begin
                    proc_path = "example.clone_vector_2_U0";
                end
                7 : begin
                    proc_path = "example.Loop_fetch_loop_proc_U0";
                end
                8 : begin
                    proc_path = "example.Loop_out_loop_proc_U0";
                end
                9 : begin
                    proc_path = "example.Loop_node_compute_lo_U0";
                end
                10 : begin
                    proc_path = "example.Loop_edge_choose_ver_U0";
                end
                11 : begin
                    proc_path = "example.Loop_edge_compute_lo_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [344:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [344:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [344:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    1: begin
                        if (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    2: begin
                        if (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    5: begin
                        if (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_example.node_attr_cpy1_V_0_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_0_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_0_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_0_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_0_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_0_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_0_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_1_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_1_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_1_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_1_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_1_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_1_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_1_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_2_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_2_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_2_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_2_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_2_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_2_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_2_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_3_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_3_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_3_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_3_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_3_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_3_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_3_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_4_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_4_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_4_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_4_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_4_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_4_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_4_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_5_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_5_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_5_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_5_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_5_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_5_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_5_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_6_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_6_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_6_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_6_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_6_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_6_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_6_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_7_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_7_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_7_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_7_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_7_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_7_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_7_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_8_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_8_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_8_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_8_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_8_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_8_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_8_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_9_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_9_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_9_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_9_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_9_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_9_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_9_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_10_s_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_10_s_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_10_s_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_10_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_10_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_10_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_10_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_10_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy1_V_10_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    9: begin
                        if (~AESL_inst_example.node_attr_cpy2_V_0_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_0_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_0_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_0_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_0_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_0_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_0_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_1_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_1_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_1_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_1_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_1_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_1_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_1_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_2_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_2_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_2_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_2_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_2_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_2_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_2_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_3_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_3_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_3_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_3_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_3_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_3_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_3_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_4_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_4_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_4_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_4_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_4_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_4_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_4_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_5_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_5_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_5_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_5_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_5_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_5_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_5_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_6_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_6_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_6_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_6_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_6_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_6_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_6_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_7_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_7_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_7_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_7_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_7_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_7_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_7_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_8_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_8_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_8_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_8_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_8_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_8_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_8_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_9_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_9_0_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_9_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_9_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_9_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_9_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_9_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_10_s_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_10_s_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_10_s_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_10_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_10_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_10_1_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_10_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_10_2_U.t_read) begin
                            chan_path = "example.node_attr_cpy2_V_10_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    0: begin
                        if (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    2: begin
                        if (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    5: begin
                        if (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    3: begin
                        if (~AESL_inst_example.edge_index_cpy1_0_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_0_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_0_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_0_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_0_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_1_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_1_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_1_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_1_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_1_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_2_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_2_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_2_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_2_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_2_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_3_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_3_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_3_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_3_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_3_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_4_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_4_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_4_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_4_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_4_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_5_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_5_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_5_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_5_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_5_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_6_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_6_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_6_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_6_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_6_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_7_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_7_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_7_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_7_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_7_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_8_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_8_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_8_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_8_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_8_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_9_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_9_0_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_9_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_9_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_9_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_10_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_10_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_10_s_U";
                            if (~AESL_inst_example.edge_index_cpy1_10_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_10_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_10_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_10_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_11_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_11_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_11_s_U";
                            if (~AESL_inst_example.edge_index_cpy1_11_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_11_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_11_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_11_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_12_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_12_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_12_s_U";
                            if (~AESL_inst_example.edge_index_cpy1_12_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_12_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_12_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_12_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy1_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_example.edge_index_cpy2_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_0_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_0_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_0_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_1_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_1_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_1_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_2_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_2_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_2_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_3_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_3_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_3_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_4_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_4_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_4_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_5_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_5_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_5_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_6_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_6_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_6_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_7_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_7_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_7_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_8_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_8_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_8_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_9_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_9_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_9_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_10_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_10_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_10_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_10_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_11_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_11_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_11_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_11_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_12_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_12_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_12_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_12_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy2_V_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    0: begin
                        if (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    1: begin
                        if (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    2: begin
                        if (~AESL_inst_example.edge_index_cpy1_0_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_0_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_0_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_0_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_0_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_1_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_1_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_1_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_1_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_1_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_2_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_2_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_2_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_2_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_2_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_3_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_3_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_3_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_3_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_3_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_4_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_4_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_4_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_4_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_4_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_5_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_5_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_5_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_5_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_5_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_6_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_6_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_6_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_6_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_6_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_7_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_7_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_7_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_7_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_7_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_8_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_8_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_8_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_8_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_8_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_9_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_9_0_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_9_0_U";
                            if (~AESL_inst_example.edge_index_cpy1_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_9_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_9_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_10_s_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_10_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_10_s_U";
                            if (~AESL_inst_example.edge_index_cpy1_10_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_10_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_10_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_10_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_11_s_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_11_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_11_s_U";
                            if (~AESL_inst_example.edge_index_cpy1_11_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_11_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_11_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_11_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_12_s_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_12_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_12_s_U";
                            if (~AESL_inst_example.edge_index_cpy1_12_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_12_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy1_12_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_12_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy1_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy1_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy1_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    7: begin
                        if (~AESL_inst_example.edge_index_cpy3_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_0_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_0_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_0_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_0_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_1_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_1_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_1_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_1_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_2_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_2_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_2_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_2_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_3_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_3_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_3_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_3_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_4_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_4_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_4_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_4_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_5_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_5_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_5_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_5_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_6_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_6_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_6_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_6_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_7_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_7_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_7_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_7_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_8_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_8_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_8_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_8_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_9_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_9_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_9_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_9_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_10_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_10_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_10_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_10_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_11_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_11_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_11_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_11_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_12_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_12_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_12_3_U.t_read) begin
                            chan_path = "example.edge_index_cpy3_V_12_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    11: begin
                        if (~AESL_inst_example.edge_index_cpy4_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_0_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_0_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_0_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_1_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_1_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_1_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_2_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_2_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_2_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_3_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_3_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_3_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_4_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_4_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_4_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_5_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_5_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_5_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_6_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_6_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_6_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_7_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_7_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_7_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_8_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_8_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_8_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_9_s_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_9_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_9_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_10_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_10_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_10_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_10_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_11_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_11_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_11_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_11_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_12_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_12_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_12_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_12_1_U.t_read) begin
                            chan_path = "example.edge_index_cpy4_V_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    1: begin
                        if (~AESL_inst_example.node_attr_cpy1_V_0_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_0_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_0_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_1_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_1_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_1_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_2_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_2_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_2_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_3_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_3_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_3_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_4_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_4_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_4_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_5_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_5_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_5_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_6_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_6_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_6_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_7_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_7_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_7_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_8_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_8_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_8_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_9_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_9_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_9_0_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_10_s_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_10_s_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_10_s_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_10_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_10_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_0_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_0_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_1_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_1_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_2_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_2_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_3_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_3_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_4_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_4_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_5_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_5_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_6_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_6_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_7_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_7_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_8_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_8_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_9_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_9_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_10_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_10_1_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_0_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_0_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_1_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_1_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_2_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_2_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_3_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_3_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_4_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_4_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_5_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_5_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_6_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_6_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_7_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_7_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_8_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_8_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_9_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_9_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy1_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_10_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy1_V_10_2_U";
                            if (~AESL_inst_example.node_attr_cpy1_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy1_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_0_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_0_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_12_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_12_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_12_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_2_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_2_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_3_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_3_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_4_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_4_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_5_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_5_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_6_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_6_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_7_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_7_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_8_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_8_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_9_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_9_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_15_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_15_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_15_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_15_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_15_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_18_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_18_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_18_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_18_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_18_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_21_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_21_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_21_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_21_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_21_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_0_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_0_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_12_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_12_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_12_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_2_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_2_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_3_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_3_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_4_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_4_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_5_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_5_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_6_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_6_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_7_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_7_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_8_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_8_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_9_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_9_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_15_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_15_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_15_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_15_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_15_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_18_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_18_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_18_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_18_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_18_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_21_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_21_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_21_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_21_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_21_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_0_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_0_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_13_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_13_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_13_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_13_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_13_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_2_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_2_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_3_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_3_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_4_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_4_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_5_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_5_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_6_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_6_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_7_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_7_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_8_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_8_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_9_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_9_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_16_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_16_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_16_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_16_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_16_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_19_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_19_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_19_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_19_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_19_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_22_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_22_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_22_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_22_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_22_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_0_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_0_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_13_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_13_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_13_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_13_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_13_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_2_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_2_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_3_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_3_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_4_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_4_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_5_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_5_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_6_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_6_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_7_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_7_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_8_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_8_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_9_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_9_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_16_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_16_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_16_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_16_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_16_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_19_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_19_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_19_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_19_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_19_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_22_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_22_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_22_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_22_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_22_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_0_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_0_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_14_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_14_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_14_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_14_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_14_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_2_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_2_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_3_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_3_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_4_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_4_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_5_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_5_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_6_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_6_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_7_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_7_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_8_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_8_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_9_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_9_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_17_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_17_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_17_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_17_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_17_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_20_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_20_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_20_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_20_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_20_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_23_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_23_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_23_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_23_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_23_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_0_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_0_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_14_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_14_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_14_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_14_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_14_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_2_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_2_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_3_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_3_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_4_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_4_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_5_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_5_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_6_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_6_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_7_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_7_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_8_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_8_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_9_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_9_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_17_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_17_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_17_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_17_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_17_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_20_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_20_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_20_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_20_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_20_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_23_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_23_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_23_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_23_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_23_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    2: begin
                        if (~AESL_inst_example.edge_index_cpy2_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_0_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_0_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_0_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_1_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_1_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_1_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_2_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_2_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_2_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_3_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_3_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_3_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_4_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_4_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_4_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_5_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_5_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_5_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_6_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_6_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_6_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_7_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_7_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_7_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_8_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_8_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_8_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_9_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_9_s_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_9_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_10_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_10_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_10_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_11_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_11_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_11_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_12_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_12_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy2_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_12_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy2_V_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy2_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy2_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    4: begin
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_0_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_0_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_0_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_0_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_0_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_0_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_12_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_12_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_12_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_12_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_13_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_13_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_13_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_13_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_13_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_13_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_13_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_13_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_13_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_13_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_14_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_14_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_14_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_14_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_14_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_14_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_14_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_14_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_14_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_14_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_2_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_2_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_2_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_2_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_2_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_2_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_3_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_3_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_3_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_3_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_3_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_3_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_4_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_4_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_4_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_4_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_4_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_4_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_5_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_5_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_5_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_5_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_5_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_5_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_6_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_6_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_6_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_6_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_6_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_6_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_7_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_7_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_7_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_7_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_7_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_7_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_8_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_8_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_8_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_8_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_8_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_8_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_9_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_9_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_9_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_9_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_9_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_9_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_15_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_15_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_15_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_15_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_15_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_15_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_15_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_15_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_15_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_15_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_16_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_16_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_16_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_16_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_16_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_16_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_16_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_16_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_16_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_16_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_17_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_17_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_17_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_17_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_17_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_17_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_17_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_17_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_17_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_17_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_18_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_18_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_18_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_18_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_18_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_18_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_18_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_18_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_18_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_18_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_19_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_19_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_19_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_19_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_19_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_19_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_19_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_19_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_19_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_19_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_20_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_20_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_20_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_20_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_20_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_20_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_20_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_20_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_20_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_20_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_21_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_21_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_21_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_21_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_21_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_21_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_21_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_21_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_21_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_21_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_22_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_22_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_22_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_22_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_22_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_22_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_22_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_22_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_22_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_22_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_23_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_23_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_23_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_23_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_23_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_23_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_23_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_23_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_23_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_23_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_example.layer7_out_0_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_0_0_V_U";
                            if (~AESL_inst_example.layer7_out_0_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_0_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_0_1_V_U";
                            if (~AESL_inst_example.layer7_out_0_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_0_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_0_2_V_U";
                            if (~AESL_inst_example.layer7_out_0_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_0_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_0_3_V_U";
                            if (~AESL_inst_example.layer7_out_0_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_1_0_V_U";
                            if (~AESL_inst_example.layer7_out_1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_1_1_V_U";
                            if (~AESL_inst_example.layer7_out_1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_1_2_V_U";
                            if (~AESL_inst_example.layer7_out_1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_1_3_V_U";
                            if (~AESL_inst_example.layer7_out_1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_2_0_V_U";
                            if (~AESL_inst_example.layer7_out_2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_2_1_V_U";
                            if (~AESL_inst_example.layer7_out_2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_2_2_V_U";
                            if (~AESL_inst_example.layer7_out_2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_2_3_V_U";
                            if (~AESL_inst_example.layer7_out_2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_3_0_V_U";
                            if (~AESL_inst_example.layer7_out_3_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_3_1_V_U";
                            if (~AESL_inst_example.layer7_out_3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_3_2_V_U";
                            if (~AESL_inst_example.layer7_out_3_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_3_3_V_U";
                            if (~AESL_inst_example.layer7_out_3_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_4_0_V_U";
                            if (~AESL_inst_example.layer7_out_4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_4_1_V_U";
                            if (~AESL_inst_example.layer7_out_4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_4_2_V_U";
                            if (~AESL_inst_example.layer7_out_4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_4_3_V_U";
                            if (~AESL_inst_example.layer7_out_4_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_5_0_V_U";
                            if (~AESL_inst_example.layer7_out_5_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_5_1_V_U";
                            if (~AESL_inst_example.layer7_out_5_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_5_2_V_U";
                            if (~AESL_inst_example.layer7_out_5_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_5_3_V_U";
                            if (~AESL_inst_example.layer7_out_5_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_6_0_V_U";
                            if (~AESL_inst_example.layer7_out_6_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_6_1_V_U";
                            if (~AESL_inst_example.layer7_out_6_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_6_2_V_U";
                            if (~AESL_inst_example.layer7_out_6_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_6_3_V_U";
                            if (~AESL_inst_example.layer7_out_6_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_7_0_V_U";
                            if (~AESL_inst_example.layer7_out_7_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_7_1_V_U";
                            if (~AESL_inst_example.layer7_out_7_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_7_2_V_U";
                            if (~AESL_inst_example.layer7_out_7_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_7_3_V_U";
                            if (~AESL_inst_example.layer7_out_7_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_8_0_V_U";
                            if (~AESL_inst_example.layer7_out_8_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_8_1_V_U";
                            if (~AESL_inst_example.layer7_out_8_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_8_2_V_U";
                            if (~AESL_inst_example.layer7_out_8_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_8_3_V_U";
                            if (~AESL_inst_example.layer7_out_8_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_9_0_V_U";
                            if (~AESL_inst_example.layer7_out_9_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_9_1_V_U";
                            if (~AESL_inst_example.layer7_out_9_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_9_2_V_U";
                            if (~AESL_inst_example.layer7_out_9_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_9_3_V_U";
                            if (~AESL_inst_example.layer7_out_9_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_10_0_V_U";
                            if (~AESL_inst_example.layer7_out_10_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_10_1_V_U";
                            if (~AESL_inst_example.layer7_out_10_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_10_2_V_U";
                            if (~AESL_inst_example.layer7_out_10_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_10_3_V_U";
                            if (~AESL_inst_example.layer7_out_10_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_11_0_V_U";
                            if (~AESL_inst_example.layer7_out_11_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_11_1_V_U";
                            if (~AESL_inst_example.layer7_out_11_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_11_2_V_U";
                            if (~AESL_inst_example.layer7_out_11_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_11_3_V_U";
                            if (~AESL_inst_example.layer7_out_11_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_0_V_U.t_read) begin
                            chan_path = "example.layer7_out_12_0_V_U";
                            if (~AESL_inst_example.layer7_out_12_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_1_V_U.t_read) begin
                            chan_path = "example.layer7_out_12_1_V_U";
                            if (~AESL_inst_example.layer7_out_12_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_2_V_U.t_read) begin
                            chan_path = "example.layer7_out_12_2_V_U";
                            if (~AESL_inst_example.layer7_out_12_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_3_V_U.t_read) begin
                            chan_path = "example.layer7_out_12_3_V_U";
                            if (~AESL_inst_example.layer7_out_12_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    0: begin
                        if (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    1: begin
                        if (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_example.layer7_out_0_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_0_0_V_U";
                            if (~AESL_inst_example.layer7_out_0_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_0_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_0_1_V_U";
                            if (~AESL_inst_example.layer7_out_0_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_0_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_0_2_V_U";
                            if (~AESL_inst_example.layer7_out_0_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_0_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_0_3_V_U";
                            if (~AESL_inst_example.layer7_out_0_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_0_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_1_0_V_U";
                            if (~AESL_inst_example.layer7_out_1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_1_1_V_U";
                            if (~AESL_inst_example.layer7_out_1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_1_2_V_U";
                            if (~AESL_inst_example.layer7_out_1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_1_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_1_3_V_U";
                            if (~AESL_inst_example.layer7_out_1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_2_0_V_U";
                            if (~AESL_inst_example.layer7_out_2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_2_1_V_U";
                            if (~AESL_inst_example.layer7_out_2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_2_2_V_U";
                            if (~AESL_inst_example.layer7_out_2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_2_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_2_3_V_U";
                            if (~AESL_inst_example.layer7_out_2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_3_0_V_U";
                            if (~AESL_inst_example.layer7_out_3_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_3_1_V_U";
                            if (~AESL_inst_example.layer7_out_3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_3_2_V_U";
                            if (~AESL_inst_example.layer7_out_3_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_3_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_3_3_V_U";
                            if (~AESL_inst_example.layer7_out_3_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_3_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_4_0_V_U";
                            if (~AESL_inst_example.layer7_out_4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_4_1_V_U";
                            if (~AESL_inst_example.layer7_out_4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_4_2_V_U";
                            if (~AESL_inst_example.layer7_out_4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_4_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_4_3_V_U";
                            if (~AESL_inst_example.layer7_out_4_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_4_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_5_0_V_U";
                            if (~AESL_inst_example.layer7_out_5_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_5_1_V_U";
                            if (~AESL_inst_example.layer7_out_5_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_5_2_V_U";
                            if (~AESL_inst_example.layer7_out_5_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_5_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_5_3_V_U";
                            if (~AESL_inst_example.layer7_out_5_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_5_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_6_0_V_U";
                            if (~AESL_inst_example.layer7_out_6_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_6_1_V_U";
                            if (~AESL_inst_example.layer7_out_6_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_6_2_V_U";
                            if (~AESL_inst_example.layer7_out_6_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_6_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_6_3_V_U";
                            if (~AESL_inst_example.layer7_out_6_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_6_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_7_0_V_U";
                            if (~AESL_inst_example.layer7_out_7_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_7_1_V_U";
                            if (~AESL_inst_example.layer7_out_7_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_7_2_V_U";
                            if (~AESL_inst_example.layer7_out_7_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_7_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_7_3_V_U";
                            if (~AESL_inst_example.layer7_out_7_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_7_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_8_0_V_U";
                            if (~AESL_inst_example.layer7_out_8_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_8_1_V_U";
                            if (~AESL_inst_example.layer7_out_8_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_8_2_V_U";
                            if (~AESL_inst_example.layer7_out_8_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_8_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_8_3_V_U";
                            if (~AESL_inst_example.layer7_out_8_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_8_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_9_0_V_U";
                            if (~AESL_inst_example.layer7_out_9_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_9_1_V_U";
                            if (~AESL_inst_example.layer7_out_9_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_9_2_V_U";
                            if (~AESL_inst_example.layer7_out_9_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_9_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_9_3_V_U";
                            if (~AESL_inst_example.layer7_out_9_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_9_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_10_0_V_U";
                            if (~AESL_inst_example.layer7_out_10_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_10_1_V_U";
                            if (~AESL_inst_example.layer7_out_10_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_10_2_V_U";
                            if (~AESL_inst_example.layer7_out_10_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_10_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_10_3_V_U";
                            if (~AESL_inst_example.layer7_out_10_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_10_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_11_0_V_U";
                            if (~AESL_inst_example.layer7_out_11_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_11_1_V_U";
                            if (~AESL_inst_example.layer7_out_11_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_11_2_V_U";
                            if (~AESL_inst_example.layer7_out_11_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_11_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_11_3_V_U";
                            if (~AESL_inst_example.layer7_out_11_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_11_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_0_V_U.i_write) begin
                            chan_path = "example.layer7_out_12_0_V_U";
                            if (~AESL_inst_example.layer7_out_12_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_1_V_U.i_write) begin
                            chan_path = "example.layer7_out_12_1_V_U";
                            if (~AESL_inst_example.layer7_out_12_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_2_V_U.i_write) begin
                            chan_path = "example.layer7_out_12_2_V_U";
                            if (~AESL_inst_example.layer7_out_12_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_12_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_3_V_U.i_write) begin
                            chan_path = "example.layer7_out_12_3_V_U";
                            if (~AESL_inst_example.layer7_out_12_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_12_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    7: begin
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_0_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_1_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_2_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_3_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_4_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_5_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_6_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_7_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_8_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_9_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_10_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_11_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_4_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_5_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_6_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_7_U.t_read) begin
                            chan_path = "example.layer7_out_cpy1_V_12_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    11: begin
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_0_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_0_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_0_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_0_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_1_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_1_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_1_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_1_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_2_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_2_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_2_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_2_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_3_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_3_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_3_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_3_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_4_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_4_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_4_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_4_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_5_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_5_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_5_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_5_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_6_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_6_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_6_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_6_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_7_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_7_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_7_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_7_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_8_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_8_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_8_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_8_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_s_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_9_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_9_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_9_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_9_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_10_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_10_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_10_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_10_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_11_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_11_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_11_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_11_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_12_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_1_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_12_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_2_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_12_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_3_U.t_read) begin
                            chan_path = "example.layer7_out_cpy2_V_12_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_example.edge_attr_aggr_0_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_0_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_1_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_2_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_3_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_4_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_5_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_6_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_7_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_8_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_9_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_10_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_11_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_1_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_2_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_3_U.t_read) begin
                            chan_path = "example.edge_attr_aggr_12_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    3: begin
                        if (~AESL_inst_example.edge_index_cpy3_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_0_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_0_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_0_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_0_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_1_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_1_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_1_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_1_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_2_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_2_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_2_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_2_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_3_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_3_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_3_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_3_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_4_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_4_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_4_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_4_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_5_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_5_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_5_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_5_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_6_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_6_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_6_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_6_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_7_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_7_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_7_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_7_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_8_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_8_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_8_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_8_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_9_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_9_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_9_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_9_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_10_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_10_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_10_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_10_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_11_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_11_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_11_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_11_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_12_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy3_V_12_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_12_3_U.i_write) begin
                            chan_path = "example.edge_index_cpy3_V_12_3_U";
                            if (~AESL_inst_example.edge_index_cpy3_V_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy3_V_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_4_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_4_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_5_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_5_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_6_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_6_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_7_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_7_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_12_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_12_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_11_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_11_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_10_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_10_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_9_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_9_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_8_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_8_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_7_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_7_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_6_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_6_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_5_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_5_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_4_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_4_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_3_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_3_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_2_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_2_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_1_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_1_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_s_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_1_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_2_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy1_V_0_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy1_V_0_3_U";
                            if (~AESL_inst_example.layer7_out_cpy1_V_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy1_V_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_example.edge_attr_aggr_0_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_0_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_0_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_1_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_2_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_1_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_3_1_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_0_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_1_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_2_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_2_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_3_2_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_0_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_0_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_0_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_0_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_1_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_1_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_1_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_1_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_2_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_2_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_2_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_2_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_3_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_3_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_3_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_3_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_4_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_4_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_4_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_4_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_5_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_5_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_5_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_5_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_6_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_6_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_6_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_6_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_7_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_7_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_7_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_7_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_8_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_8_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_8_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_8_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_9_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_9_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_9_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_9_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_10_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_10_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_10_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_10_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_11_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_11_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_11_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_11_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_0_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_1_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_2_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_attr_aggr_12_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_3_U.i_write) begin
                            chan_path = "example.edge_attr_aggr_12_3_3_U";
                            if (~AESL_inst_example.edge_attr_aggr_12_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_attr_aggr_12_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    9: begin
                        if (~AESL_inst_example.layer9_out_1_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_1_0_V_U";
                            if (~AESL_inst_example.layer9_out_1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_2_0_V_U";
                            if (~AESL_inst_example.layer9_out_2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_3_0_V_U";
                            if (~AESL_inst_example.layer9_out_3_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_4_0_V_U";
                            if (~AESL_inst_example.layer9_out_4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_5_0_V_U";
                            if (~AESL_inst_example.layer9_out_5_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_6_0_V_U";
                            if (~AESL_inst_example.layer9_out_6_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_7_0_V_U";
                            if (~AESL_inst_example.layer9_out_7_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_8_0_V_U";
                            if (~AESL_inst_example.layer9_out_8_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_9_0_V_U";
                            if (~AESL_inst_example.layer9_out_9_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_0_V_U.t_read) begin
                            chan_path = "example.layer9_out_10_0_V_U";
                            if (~AESL_inst_example.layer9_out_10_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_1_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_1_1_V_U";
                            if (~AESL_inst_example.layer9_out_1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_2_1_V_U";
                            if (~AESL_inst_example.layer9_out_2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_3_1_V_U";
                            if (~AESL_inst_example.layer9_out_3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_4_1_V_U";
                            if (~AESL_inst_example.layer9_out_4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_5_1_V_U";
                            if (~AESL_inst_example.layer9_out_5_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_6_1_V_U";
                            if (~AESL_inst_example.layer9_out_6_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_7_1_V_U";
                            if (~AESL_inst_example.layer9_out_7_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_8_1_V_U";
                            if (~AESL_inst_example.layer9_out_8_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_9_1_V_U";
                            if (~AESL_inst_example.layer9_out_9_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_1_V_U.t_read) begin
                            chan_path = "example.layer9_out_10_1_V_U";
                            if (~AESL_inst_example.layer9_out_10_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_1_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_1_2_V_U";
                            if (~AESL_inst_example.layer9_out_1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_2_2_V_U";
                            if (~AESL_inst_example.layer9_out_2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_3_2_V_U";
                            if (~AESL_inst_example.layer9_out_3_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_4_2_V_U";
                            if (~AESL_inst_example.layer9_out_4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_5_2_V_U";
                            if (~AESL_inst_example.layer9_out_5_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_6_2_V_U";
                            if (~AESL_inst_example.layer9_out_6_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_7_2_V_U";
                            if (~AESL_inst_example.layer9_out_7_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_8_2_V_U";
                            if (~AESL_inst_example.layer9_out_8_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_9_2_V_U";
                            if (~AESL_inst_example.layer9_out_9_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_2_V_U.t_read) begin
                            chan_path = "example.layer9_out_10_2_V_U";
                            if (~AESL_inst_example.layer9_out_10_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_1_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_1_3_V_U";
                            if (~AESL_inst_example.layer9_out_1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_2_3_V_U";
                            if (~AESL_inst_example.layer9_out_2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_3_3_V_U";
                            if (~AESL_inst_example.layer9_out_3_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_4_3_V_U";
                            if (~AESL_inst_example.layer9_out_4_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_5_3_V_U";
                            if (~AESL_inst_example.layer9_out_5_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_6_3_V_U";
                            if (~AESL_inst_example.layer9_out_6_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_7_3_V_U";
                            if (~AESL_inst_example.layer9_out_7_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_8_3_V_U";
                            if (~AESL_inst_example.layer9_out_8_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_9_3_V_U";
                            if (~AESL_inst_example.layer9_out_9_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_3_V_U.t_read) begin
                            chan_path = "example.layer9_out_10_3_V_U";
                            if (~AESL_inst_example.layer9_out_10_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    1: begin
                        if (~AESL_inst_example.node_attr_cpy2_V_0_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_0_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_0_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_0_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_0_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_0_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_0_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_0_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_0_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_1_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_1_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_1_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_1_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_1_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_1_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_1_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_1_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_1_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_2_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_2_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_2_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_2_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_2_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_2_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_2_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_2_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_2_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_3_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_3_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_3_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_3_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_3_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_3_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_3_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_3_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_3_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_4_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_4_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_4_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_4_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_4_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_4_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_4_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_4_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_4_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_5_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_5_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_5_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_5_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_5_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_5_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_5_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_5_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_5_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_6_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_6_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_6_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_6_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_6_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_6_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_6_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_6_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_6_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_7_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_7_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_7_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_7_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_7_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_7_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_7_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_7_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_7_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_8_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_8_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_8_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_8_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_8_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_8_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_8_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_8_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_8_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_9_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_9_0_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_9_0_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_9_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_9_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_9_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_9_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_9_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_9_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_10_s_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_10_s_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_10_s_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_10_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_10_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_10_1_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_10_1_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_cpy2_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_10_2_U.i_write) begin
                            chan_path = "example.node_attr_cpy2_V_10_2_U";
                            if (~AESL_inst_example.node_attr_cpy2_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_cpy2_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_example.layer10_out_0_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_0_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_0_0_V_U";
                            if (~AESL_inst_example.layer10_out_0_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_0_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_0_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_0_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_0_1_V_U";
                            if (~AESL_inst_example.layer10_out_0_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_0_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_0_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_0_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_0_2_V_U";
                            if (~AESL_inst_example.layer10_out_0_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_0_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_1_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_1_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_1_0_V_U";
                            if (~AESL_inst_example.layer10_out_1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_1_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_1_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_1_1_V_U";
                            if (~AESL_inst_example.layer10_out_1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_1_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_1_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_1_2_V_U";
                            if (~AESL_inst_example.layer10_out_1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_2_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_2_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_2_0_V_U";
                            if (~AESL_inst_example.layer10_out_2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_2_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_2_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_2_1_V_U";
                            if (~AESL_inst_example.layer10_out_2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_2_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_2_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_2_2_V_U";
                            if (~AESL_inst_example.layer10_out_2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_3_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_3_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_3_0_V_U";
                            if (~AESL_inst_example.layer10_out_3_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_3_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_3_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_3_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_3_1_V_U";
                            if (~AESL_inst_example.layer10_out_3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_3_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_3_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_3_2_V_U";
                            if (~AESL_inst_example.layer10_out_3_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_3_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_4_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_4_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_4_0_V_U";
                            if (~AESL_inst_example.layer10_out_4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_4_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_4_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_4_1_V_U";
                            if (~AESL_inst_example.layer10_out_4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_4_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_4_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_4_2_V_U";
                            if (~AESL_inst_example.layer10_out_4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_5_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_5_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_5_0_V_U";
                            if (~AESL_inst_example.layer10_out_5_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_5_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_5_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_5_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_5_1_V_U";
                            if (~AESL_inst_example.layer10_out_5_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_5_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_5_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_5_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_5_2_V_U";
                            if (~AESL_inst_example.layer10_out_5_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_5_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_6_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_6_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_6_0_V_U";
                            if (~AESL_inst_example.layer10_out_6_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_6_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_6_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_6_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_6_1_V_U";
                            if (~AESL_inst_example.layer10_out_6_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_6_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_6_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_6_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_6_2_V_U";
                            if (~AESL_inst_example.layer10_out_6_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_6_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_7_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_7_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_7_0_V_U";
                            if (~AESL_inst_example.layer10_out_7_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_7_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_7_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_7_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_7_1_V_U";
                            if (~AESL_inst_example.layer10_out_7_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_7_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_7_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_7_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_7_2_V_U";
                            if (~AESL_inst_example.layer10_out_7_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_7_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_8_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_8_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_8_0_V_U";
                            if (~AESL_inst_example.layer10_out_8_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_8_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_8_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_8_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_8_1_V_U";
                            if (~AESL_inst_example.layer10_out_8_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_8_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_8_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_8_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_8_2_V_U";
                            if (~AESL_inst_example.layer10_out_8_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_8_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_9_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_9_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_9_0_V_U";
                            if (~AESL_inst_example.layer10_out_9_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_9_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_9_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_9_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_9_1_V_U";
                            if (~AESL_inst_example.layer10_out_9_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_9_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_9_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_9_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_9_2_V_U";
                            if (~AESL_inst_example.layer10_out_9_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_9_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_10_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_10_0_V_U.t_read) begin
                            chan_path = "example.layer10_out_10_0_V_U";
                            if (~AESL_inst_example.layer10_out_10_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_10_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_10_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_10_1_V_U.t_read) begin
                            chan_path = "example.layer10_out_10_1_V_U";
                            if (~AESL_inst_example.layer10_out_10_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_10_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_10_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_10_2_V_U.t_read) begin
                            chan_path = "example.layer10_out_10_2_V_U";
                            if (~AESL_inst_example.layer10_out_10_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_10_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    8: begin
                        if (~AESL_inst_example.layer9_out_1_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_1_0_V_U";
                            if (~AESL_inst_example.layer9_out_1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_1_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_1_1_V_U";
                            if (~AESL_inst_example.layer9_out_1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_1_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_1_2_V_U";
                            if (~AESL_inst_example.layer9_out_1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_1_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_1_3_V_U";
                            if (~AESL_inst_example.layer9_out_1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_2_0_V_U";
                            if (~AESL_inst_example.layer9_out_2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_2_1_V_U";
                            if (~AESL_inst_example.layer9_out_2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_2_2_V_U";
                            if (~AESL_inst_example.layer9_out_2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_2_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_2_3_V_U";
                            if (~AESL_inst_example.layer9_out_2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_3_0_V_U";
                            if (~AESL_inst_example.layer9_out_3_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_3_1_V_U";
                            if (~AESL_inst_example.layer9_out_3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_3_2_V_U";
                            if (~AESL_inst_example.layer9_out_3_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_3_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_3_3_V_U";
                            if (~AESL_inst_example.layer9_out_3_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_3_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_4_0_V_U";
                            if (~AESL_inst_example.layer9_out_4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_4_1_V_U";
                            if (~AESL_inst_example.layer9_out_4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_4_2_V_U";
                            if (~AESL_inst_example.layer9_out_4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_4_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_4_3_V_U";
                            if (~AESL_inst_example.layer9_out_4_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_4_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_5_0_V_U";
                            if (~AESL_inst_example.layer9_out_5_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_5_1_V_U";
                            if (~AESL_inst_example.layer9_out_5_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_5_2_V_U";
                            if (~AESL_inst_example.layer9_out_5_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_5_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_5_3_V_U";
                            if (~AESL_inst_example.layer9_out_5_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_5_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_6_0_V_U";
                            if (~AESL_inst_example.layer9_out_6_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_6_1_V_U";
                            if (~AESL_inst_example.layer9_out_6_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_6_2_V_U";
                            if (~AESL_inst_example.layer9_out_6_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_6_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_6_3_V_U";
                            if (~AESL_inst_example.layer9_out_6_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_6_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_7_0_V_U";
                            if (~AESL_inst_example.layer9_out_7_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_7_1_V_U";
                            if (~AESL_inst_example.layer9_out_7_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_7_2_V_U";
                            if (~AESL_inst_example.layer9_out_7_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_7_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_7_3_V_U";
                            if (~AESL_inst_example.layer9_out_7_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_7_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_8_0_V_U";
                            if (~AESL_inst_example.layer9_out_8_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_8_1_V_U";
                            if (~AESL_inst_example.layer9_out_8_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_8_2_V_U";
                            if (~AESL_inst_example.layer9_out_8_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_8_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_8_3_V_U";
                            if (~AESL_inst_example.layer9_out_8_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_8_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_9_0_V_U";
                            if (~AESL_inst_example.layer9_out_9_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_9_1_V_U";
                            if (~AESL_inst_example.layer9_out_9_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_9_2_V_U";
                            if (~AESL_inst_example.layer9_out_9_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_9_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_9_3_V_U";
                            if (~AESL_inst_example.layer9_out_9_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_9_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_0_V_U.i_write) begin
                            chan_path = "example.layer9_out_10_0_V_U";
                            if (~AESL_inst_example.layer9_out_10_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_1_V_U.i_write) begin
                            chan_path = "example.layer9_out_10_1_V_U";
                            if (~AESL_inst_example.layer9_out_10_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_2_V_U.i_write) begin
                            chan_path = "example.layer9_out_10_2_V_U";
                            if (~AESL_inst_example.layer9_out_10_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer9_out_10_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_3_V_U.i_write) begin
                            chan_path = "example.layer9_out_10_3_V_U";
                            if (~AESL_inst_example.layer9_out_10_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer9_out_10_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    9: begin
                        if (~AESL_inst_example.layer10_out_0_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_0_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_0_0_V_U";
                            if (~AESL_inst_example.layer10_out_0_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_0_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_1_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_1_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_1_0_V_U";
                            if (~AESL_inst_example.layer10_out_1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_2_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_2_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_2_0_V_U";
                            if (~AESL_inst_example.layer10_out_2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_3_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_3_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_3_0_V_U";
                            if (~AESL_inst_example.layer10_out_3_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_3_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_4_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_4_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_4_0_V_U";
                            if (~AESL_inst_example.layer10_out_4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_5_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_5_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_5_0_V_U";
                            if (~AESL_inst_example.layer10_out_5_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_5_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_6_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_6_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_6_0_V_U";
                            if (~AESL_inst_example.layer10_out_6_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_6_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_7_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_7_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_7_0_V_U";
                            if (~AESL_inst_example.layer10_out_7_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_7_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_8_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_8_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_8_0_V_U";
                            if (~AESL_inst_example.layer10_out_8_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_8_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_9_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_9_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_9_0_V_U";
                            if (~AESL_inst_example.layer10_out_9_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_9_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_10_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_10_0_V_U.i_write) begin
                            chan_path = "example.layer10_out_10_0_V_U";
                            if (~AESL_inst_example.layer10_out_10_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_10_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_0_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_0_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_0_1_V_U";
                            if (~AESL_inst_example.layer10_out_0_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_0_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_1_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_1_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_1_1_V_U";
                            if (~AESL_inst_example.layer10_out_1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_2_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_2_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_2_1_V_U";
                            if (~AESL_inst_example.layer10_out_2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_3_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_3_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_3_1_V_U";
                            if (~AESL_inst_example.layer10_out_3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_4_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_4_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_4_1_V_U";
                            if (~AESL_inst_example.layer10_out_4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_5_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_5_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_5_1_V_U";
                            if (~AESL_inst_example.layer10_out_5_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_5_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_6_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_6_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_6_1_V_U";
                            if (~AESL_inst_example.layer10_out_6_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_6_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_7_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_7_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_7_1_V_U";
                            if (~AESL_inst_example.layer10_out_7_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_7_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_8_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_8_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_8_1_V_U";
                            if (~AESL_inst_example.layer10_out_8_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_8_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_9_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_9_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_9_1_V_U";
                            if (~AESL_inst_example.layer10_out_9_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_9_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_10_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_10_1_V_U.i_write) begin
                            chan_path = "example.layer10_out_10_1_V_U";
                            if (~AESL_inst_example.layer10_out_10_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_10_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_0_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_0_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_0_2_V_U";
                            if (~AESL_inst_example.layer10_out_0_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_0_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_1_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_1_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_1_2_V_U";
                            if (~AESL_inst_example.layer10_out_1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_2_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_2_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_2_2_V_U";
                            if (~AESL_inst_example.layer10_out_2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_3_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_3_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_3_2_V_U";
                            if (~AESL_inst_example.layer10_out_3_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_3_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_4_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_4_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_4_2_V_U";
                            if (~AESL_inst_example.layer10_out_4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_5_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_5_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_5_2_V_U";
                            if (~AESL_inst_example.layer10_out_5_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_5_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_6_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_6_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_6_2_V_U";
                            if (~AESL_inst_example.layer10_out_6_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_6_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_7_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_7_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_7_2_V_U";
                            if (~AESL_inst_example.layer10_out_7_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_7_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_8_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_8_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_8_2_V_U";
                            if (~AESL_inst_example.layer10_out_8_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_8_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_9_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_9_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_9_2_V_U";
                            if (~AESL_inst_example.layer10_out_9_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_9_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer10_out_10_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_10_2_V_U.i_write) begin
                            chan_path = "example.layer10_out_10_2_V_U";
                            if (~AESL_inst_example.layer10_out_10_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer10_out_10_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    11: begin
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_0_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_0_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_6_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_6_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_7_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_7_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_8_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_8_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_9_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_9_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_6_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_6_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_9_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_9_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_0_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_0_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_6_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_6_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_7_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_7_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_8_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_8_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_9_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_9_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_3_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_6_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_6_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_9_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_9_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_0_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_0_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_2_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_2_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_3_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_3_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_4_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_4_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_5_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_5_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_6_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_6_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_7_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_7_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_8_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_8_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_9_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_9_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_7_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_7_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_10_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_10_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_10_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_0_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_0_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_2_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_2_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_3_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_3_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_4_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_4_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_5_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_5_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_6_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_6_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_7_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_7_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_8_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_8_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_9_1_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_9_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_4_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_7_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_7_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_10_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_10_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_10_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_0_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_0_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_2_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_2_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_3_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_3_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_4_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_4_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_5_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_5_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_6_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_6_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_7_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_7_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_8_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_8_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_9_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_9_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_8_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_8_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_11_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_11_U.t_read) begin
                            chan_path = "example.node_attr_1D_s_mat_1_11_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_0_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_0_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_2_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_2_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_3_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_3_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_4_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_4_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_5_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_5_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_6_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_6_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_7_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_7_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_8_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_8_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_9_2_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_9_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_5_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_8_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_8_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_11_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_11_U.t_read) begin
                            chan_path = "example.node_attr_1D_r_mat_1_11_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    6: begin
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_0_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_0_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_0_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_0_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_0_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_0_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_0_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_1_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_1_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_1_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_1_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_1_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_2_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_2_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_2_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_2_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_2_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_2_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_2_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_3_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_3_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_3_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_3_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_3_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_3_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_3_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_4_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_4_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_4_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_4_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_4_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_4_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_4_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_5_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_5_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_5_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_5_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_5_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_5_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_5_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_6_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_6_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_6_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_6_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_6_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_6_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_6_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_7_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_7_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_7_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_7_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_7_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_7_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_7_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_8_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_8_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_8_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_8_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_8_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_8_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_8_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_s_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_9_s_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_9_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_9_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_9_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_9_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_9_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_9_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_10_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_10_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_10_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_10_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_10_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_10_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_10_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_11_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_11_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_11_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_11_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_11_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_11_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_11_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_12_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_1_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_12_1_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_2_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_12_2_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.layer7_out_cpy2_V_12_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_3_U.i_write) begin
                            chan_path = "example.layer7_out_cpy2_V_12_3_U";
                            if (~AESL_inst_example.layer7_out_cpy2_V_12_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.layer7_out_cpy2_V_12_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    3: begin
                        if (~AESL_inst_example.edge_index_cpy4_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_0_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_0_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_0_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_0_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_0_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_0_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_1_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_1_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_1_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_1_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_1_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_1_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_2_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_2_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_2_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_2_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_2_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_2_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_3_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_3_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_3_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_3_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_3_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_3_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_4_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_4_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_4_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_4_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_4_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_4_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_5_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_5_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_5_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_5_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_5_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_5_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_6_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_6_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_6_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_6_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_6_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_6_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_7_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_7_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_7_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_7_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_7_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_7_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_8_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_8_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_8_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_8_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_8_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_8_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_9_s_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_9_s_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_9_s_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_9_s_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_9_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_9_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_10_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_10_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_10_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_10_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_10_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_10_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_11_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_11_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_11_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_11_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_11_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_11_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_12_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_12_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_12_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_12_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.edge_index_cpy4_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_12_1_U.i_write) begin
                            chan_path = "example.edge_index_cpy4_V_12_1_U";
                            if (~AESL_inst_example.edge_index_cpy4_V_12_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.edge_index_cpy4_V_12_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_0_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_0_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_0_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_0_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_0_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_0_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_0_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_0_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_2_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_2_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_2_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_2_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_2_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_2_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_3_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_3_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_3_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_3_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_3_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_3_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_4_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_4_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_4_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_4_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_4_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_4_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_5_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_5_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_5_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_5_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_5_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_5_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_6_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_6_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_6_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_6_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_6_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_6_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_6_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_6_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_7_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_7_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_7_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_7_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_7_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_7_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_7_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_7_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_8_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_8_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_8_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_8_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_8_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_8_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_8_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_8_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_9_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_9_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_9_1_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_1_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_9_1_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_1_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_1_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_9_2_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_2_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_9_2_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_9_2_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_9_2_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_3_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_3_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_3_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_3_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_3_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_4_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_4_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_4_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_4_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_4_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_5_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_5_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_5_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_5_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_5_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_6_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_6_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_6_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_6_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_6_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_6_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_7_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_7_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_7_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_7_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_7_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_7_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_8_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_8_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_8_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_8_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_8_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_8_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_9_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_9_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_9_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_9_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_9_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_9_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_10_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_10_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_10_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_10_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_10_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_10_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_s_mat_1_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_11_U.i_write) begin
                            chan_path = "example.node_attr_1D_s_mat_1_11_U";
                            if (~AESL_inst_example.node_attr_1D_s_mat_1_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_s_mat_1_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_example.node_attr_1D_r_mat_1_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_11_U.i_write) begin
                            chan_path = "example.node_attr_1D_r_mat_1_11_U";
                            if (~AESL_inst_example.node_attr_1D_r_mat_1_11_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_example.node_attr_1D_r_mat_1_11_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        wait (reset == 1);
        cycle_id = 1;
        while (1) begin
            @ (negedge clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end(cycle_id - 1);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
endmodule
