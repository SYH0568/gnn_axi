`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input reset,
    input clock);

    wire [2:0] proc_dep_vld_vec_0;
    reg [2:0] proc_dep_vld_vec_0_reg;
    wire [2:0] in_chan_dep_vld_vec_0;
    wire [35:0] in_chan_dep_data_vec_0;
    wire [2:0] token_in_vec_0;
    wire [2:0] out_chan_dep_vld_vec_0;
    wire [11:0] out_chan_dep_data_0;
    wire [2:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [11:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [11:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_5_0;
    wire [11:0] dep_chan_data_5_0;
    wire token_5_0;
    wire [4:0] proc_dep_vld_vec_1;
    reg [4:0] proc_dep_vld_vec_1_reg;
    wire [4:0] in_chan_dep_vld_vec_1;
    wire [59:0] in_chan_dep_data_vec_1;
    wire [4:0] token_in_vec_1;
    wire [4:0] out_chan_dep_vld_vec_1;
    wire [11:0] out_chan_dep_data_1;
    wire [4:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [11:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [11:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_4_1;
    wire [11:0] dep_chan_data_4_1;
    wire token_4_1;
    wire dep_chan_vld_5_1;
    wire [11:0] dep_chan_data_5_1;
    wire token_5_1;
    wire dep_chan_vld_9_1;
    wire [11:0] dep_chan_data_9_1;
    wire token_9_1;
    wire [3:0] proc_dep_vld_vec_2;
    reg [3:0] proc_dep_vld_vec_2_reg;
    wire [3:0] in_chan_dep_vld_vec_2;
    wire [47:0] in_chan_dep_data_vec_2;
    wire [3:0] token_in_vec_2;
    wire [3:0] out_chan_dep_vld_vec_2;
    wire [11:0] out_chan_dep_data_2;
    wire [3:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [11:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [11:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_3_2;
    wire [11:0] dep_chan_data_3_2;
    wire token_3_2;
    wire dep_chan_vld_5_2;
    wire [11:0] dep_chan_data_5_2;
    wire token_5_2;
    wire [2:0] proc_dep_vld_vec_3;
    reg [2:0] proc_dep_vld_vec_3_reg;
    wire [2:0] in_chan_dep_vld_vec_3;
    wire [35:0] in_chan_dep_data_vec_3;
    wire [2:0] token_in_vec_3;
    wire [2:0] out_chan_dep_vld_vec_3;
    wire [11:0] out_chan_dep_data_3;
    wire [2:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_2_3;
    wire [11:0] dep_chan_data_2_3;
    wire token_2_3;
    wire dep_chan_vld_7_3;
    wire [11:0] dep_chan_data_7_3;
    wire token_7_3;
    wire dep_chan_vld_11_3;
    wire [11:0] dep_chan_data_11_3;
    wire token_11_3;
    wire [1:0] proc_dep_vld_vec_4;
    reg [1:0] proc_dep_vld_vec_4_reg;
    wire [1:0] in_chan_dep_vld_vec_4;
    wire [23:0] in_chan_dep_data_vec_4;
    wire [1:0] token_in_vec_4;
    wire [1:0] out_chan_dep_vld_vec_4;
    wire [11:0] out_chan_dep_data_4;
    wire [1:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_1_4;
    wire [11:0] dep_chan_data_1_4;
    wire token_1_4;
    wire dep_chan_vld_5_4;
    wire [11:0] dep_chan_data_5_4;
    wire token_5_4;
    wire [4:0] proc_dep_vld_vec_5;
    reg [4:0] proc_dep_vld_vec_5_reg;
    wire [4:0] in_chan_dep_vld_vec_5;
    wire [59:0] in_chan_dep_data_vec_5;
    wire [4:0] token_in_vec_5;
    wire [4:0] out_chan_dep_vld_vec_5;
    wire [11:0] out_chan_dep_data_5;
    wire [4:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_0_5;
    wire [11:0] dep_chan_data_0_5;
    wire token_0_5;
    wire dep_chan_vld_1_5;
    wire [11:0] dep_chan_data_1_5;
    wire token_1_5;
    wire dep_chan_vld_2_5;
    wire [11:0] dep_chan_data_2_5;
    wire token_2_5;
    wire dep_chan_vld_4_5;
    wire [11:0] dep_chan_data_4_5;
    wire token_4_5;
    wire dep_chan_vld_6_5;
    wire [11:0] dep_chan_data_6_5;
    wire token_6_5;
    wire [2:0] proc_dep_vld_vec_6;
    reg [2:0] proc_dep_vld_vec_6_reg;
    wire [2:0] in_chan_dep_vld_vec_6;
    wire [35:0] in_chan_dep_data_vec_6;
    wire [2:0] token_in_vec_6;
    wire [2:0] out_chan_dep_vld_vec_6;
    wire [11:0] out_chan_dep_data_6;
    wire [2:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_5_6;
    wire [11:0] dep_chan_data_5_6;
    wire token_5_6;
    wire dep_chan_vld_7_6;
    wire [11:0] dep_chan_data_7_6;
    wire token_7_6;
    wire dep_chan_vld_11_6;
    wire [11:0] dep_chan_data_11_6;
    wire token_11_6;
    wire [2:0] proc_dep_vld_vec_7;
    reg [2:0] proc_dep_vld_vec_7_reg;
    wire [2:0] in_chan_dep_vld_vec_7;
    wire [35:0] in_chan_dep_data_vec_7;
    wire [2:0] token_in_vec_7;
    wire [2:0] out_chan_dep_vld_vec_7;
    wire [11:0] out_chan_dep_data_7;
    wire [2:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_3_7;
    wire [11:0] dep_chan_data_3_7;
    wire token_3_7;
    wire dep_chan_vld_6_7;
    wire [11:0] dep_chan_data_6_7;
    wire token_6_7;
    wire dep_chan_vld_8_7;
    wire [11:0] dep_chan_data_8_7;
    wire token_8_7;
    wire [1:0] proc_dep_vld_vec_8;
    reg [1:0] proc_dep_vld_vec_8_reg;
    wire [1:0] in_chan_dep_vld_vec_8;
    wire [23:0] in_chan_dep_data_vec_8;
    wire [1:0] token_in_vec_8;
    wire [1:0] out_chan_dep_vld_vec_8;
    wire [11:0] out_chan_dep_data_8;
    wire [1:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_7_8;
    wire [11:0] dep_chan_data_7_8;
    wire token_7_8;
    wire dep_chan_vld_9_8;
    wire [11:0] dep_chan_data_9_8;
    wire token_9_8;
    wire [2:0] proc_dep_vld_vec_9;
    reg [2:0] proc_dep_vld_vec_9_reg;
    wire [2:0] in_chan_dep_vld_vec_9;
    wire [35:0] in_chan_dep_data_vec_9;
    wire [2:0] token_in_vec_9;
    wire [2:0] out_chan_dep_vld_vec_9;
    wire [11:0] out_chan_dep_data_9;
    wire [2:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_1_9;
    wire [11:0] dep_chan_data_1_9;
    wire token_1_9;
    wire dep_chan_vld_8_9;
    wire [11:0] dep_chan_data_8_9;
    wire token_8_9;
    wire dep_chan_vld_10_9;
    wire [11:0] dep_chan_data_10_9;
    wire token_10_9;
    wire [1:0] proc_dep_vld_vec_10;
    reg [1:0] proc_dep_vld_vec_10_reg;
    wire [1:0] in_chan_dep_vld_vec_10;
    wire [23:0] in_chan_dep_data_vec_10;
    wire [1:0] token_in_vec_10;
    wire [1:0] out_chan_dep_vld_vec_10;
    wire [11:0] out_chan_dep_data_10;
    wire [1:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_9_10;
    wire [11:0] dep_chan_data_9_10;
    wire token_9_10;
    wire dep_chan_vld_11_10;
    wire [11:0] dep_chan_data_11_10;
    wire token_11_10;
    wire [2:0] proc_dep_vld_vec_11;
    reg [2:0] proc_dep_vld_vec_11_reg;
    wire [2:0] in_chan_dep_vld_vec_11;
    wire [35:0] in_chan_dep_data_vec_11;
    wire [2:0] token_in_vec_11;
    wire [2:0] out_chan_dep_vld_vec_11;
    wire [11:0] out_chan_dep_data_11;
    wire [2:0] token_out_vec_11;
    wire dl_detect_out_11;
    wire dep_chan_vld_3_11;
    wire [11:0] dep_chan_data_3_11;
    wire token_3_11;
    wire dep_chan_vld_6_11;
    wire [11:0] dep_chan_data_6_11;
    wire token_6_11;
    wire dep_chan_vld_10_11;
    wire [11:0] dep_chan_data_10_11;
    wire token_10_11;
    wire [11:0] dl_in_vec;
    wire dl_detect_out;
    wire [11:0] origin;
    wire token_clear;

    reg ap_done_reg_0;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_example.clone_vector_3_U0.ap_done;
        end
    end

    reg ap_done_reg_1;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_example.clone_vector_1_U0.ap_done;
        end
    end

    reg ap_done_reg_2;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_2 <= 'b0;
        end
        else begin
            ap_done_reg_2 <= AESL_inst_example.clone_vector_U0.ap_done;
        end
    end

    reg ap_done_reg_3;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_3 <= 'b0;
        end
        else begin
            ap_done_reg_3 <= AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done;
        end
    end

    reg ap_done_reg_4;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_4 <= 'b0;
        end
        else begin
            ap_done_reg_4 <= AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done;
        end
    end

    reg ap_done_reg_5;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_5 <= 'b0;
        end
        else begin
            ap_done_reg_5 <= AESL_inst_example.clone_vector_2_U0.ap_done;
        end
    end

    reg ap_done_reg_6;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_6 <= 'b0;
        end
        else begin
            ap_done_reg_6 <= AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done;
        end
    end

    reg ap_done_reg_7;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_7 <= 'b0;
        end
        else begin
            ap_done_reg_7 <= AESL_inst_example.Loop_out_loop_proc_U0.ap_done;
        end
    end

    reg ap_done_reg_8;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_8 <= 'b0;
        end
        else begin
            ap_done_reg_8 <= AESL_inst_example.Loop_node_compute_lo_U0.ap_done;
        end
    end

    reg ap_done_reg_9;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_9 <= 'b0;
        end
        else begin
            ap_done_reg_9 <= AESL_inst_example.Loop_edge_choose_ver_U0.ap_done;
        end
    end

    reg ap_done_reg_10;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_10 <= 'b0;
        end
        else begin
            ap_done_reg_10 <= AESL_inst_example.Loop_edge_compute_lo_U0.ap_done;
        end
    end

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Block_proc_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Block_proc_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Block_proc_U0$ap_idle <= AESL_inst_example.Block_proc_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Block_proc_U0
    AESL_deadlock_detect_unit #(12, 0, 3, 3) AESL_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (((AESL_inst_example.Block_proc_U0_ap_ready_count[0]) & AESL_inst_example.Block_proc_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[11 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[23 : 12] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_5_0;
    assign in_chan_dep_data_vec_0[35 : 24] = dep_chan_data_5_0;
    assign token_in_vec_0[2] = token_5_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[1];
    assign dep_chan_vld_0_5 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_5 = out_chan_dep_data_0;
    assign token_0_5 = token_out_vec_0[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$clone_vector_3_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$clone_vector_3_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$clone_vector_3_U0$ap_idle <= AESL_inst_example.clone_vector_3_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.clone_vector_3_U0
    AESL_deadlock_detect_unit #(12, 1, 5, 5) AESL_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (~AESL_inst_example.node_attr_cpy1_V_0_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_0_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_0_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_0_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_1_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_1_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_1_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_1_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_2_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_2_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_2_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_2_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_3_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_3_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_3_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_3_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_4_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_4_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_4_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_4_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_5_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_5_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_5_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_5_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_6_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_6_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_6_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_6_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_7_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_7_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_7_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_7_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_8_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_8_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_8_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_8_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_9_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_9_0_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_9_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_9_2_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_10_s_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_10_s_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_10_1_U.t_read | ~AESL_inst_example.node_attr_cpy1_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy1_V_10_2_U.t_read);
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (~AESL_inst_example.node_attr_cpy2_V_0_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_0_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_0_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_0_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_1_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_1_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_1_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_1_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_2_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_2_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_2_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_2_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_3_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_3_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_3_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_3_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_4_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_4_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_4_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_4_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_5_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_5_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_5_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_5_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_6_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_6_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_6_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_6_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_7_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_7_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_7_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_7_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_8_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_8_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_8_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_8_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_9_0_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_9_0_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_9_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_9_2_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_10_s_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_10_s_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_10_1_U.t_read | ~AESL_inst_example.node_attr_cpy2_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_3_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_example.node_attr_cpy2_V_10_2_U.t_read);
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_1[4] = dl_detect_out ? proc_dep_vld_vec_1_reg[4] : (((AESL_inst_example.clone_vector_3_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_3_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[11 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[23 : 12] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_4_1;
    assign in_chan_dep_data_vec_1[35 : 24] = dep_chan_data_4_1;
    assign token_in_vec_1[2] = token_4_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_5_1;
    assign in_chan_dep_data_vec_1[47 : 36] = dep_chan_data_5_1;
    assign token_in_vec_1[3] = token_5_1;
    assign in_chan_dep_vld_vec_1[4] = dep_chan_vld_9_1;
    assign in_chan_dep_data_vec_1[59 : 48] = dep_chan_data_9_1;
    assign token_in_vec_1[4] = token_9_1;
    assign dep_chan_vld_1_4 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_4 = out_chan_dep_data_1;
    assign token_1_4 = token_out_vec_1[0];
    assign dep_chan_vld_1_9 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_9 = out_chan_dep_data_1;
    assign token_1_9 = token_out_vec_1[1];
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[2];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[3];
    assign dep_chan_vld_1_5 = out_chan_dep_vld_vec_1[4];
    assign dep_chan_data_1_5 = out_chan_dep_data_1;
    assign token_1_5 = token_out_vec_1[4];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$clone_vector_1_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$clone_vector_1_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$clone_vector_1_U0$ap_idle <= AESL_inst_example.clone_vector_1_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.clone_vector_1_U0
    AESL_deadlock_detect_unit #(12, 2, 4, 4) AESL_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (~AESL_inst_example.edge_index_cpy1_0_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_0_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_0_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_0_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_1_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_1_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_1_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_1_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_2_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_2_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_2_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_2_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_3_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_3_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_3_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_3_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_4_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_4_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_4_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_4_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_5_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_5_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_5_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_5_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_6_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_6_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_6_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_6_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_7_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_7_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_7_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_7_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_8_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_8_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_8_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_8_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_9_0_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_9_0_U.t_read | ~AESL_inst_example.edge_index_cpy1_9_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_9_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_10_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_10_s_U.t_read | ~AESL_inst_example.edge_index_cpy1_10_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_10_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_11_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_11_s_U.t_read | ~AESL_inst_example.edge_index_cpy1_11_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_11_1_U.t_read | ~AESL_inst_example.edge_index_cpy1_12_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_12_s_U.t_read | ~AESL_inst_example.edge_index_cpy1_12_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy1_12_1_U.t_read);
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (~AESL_inst_example.edge_index_cpy2_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_0_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_0_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_1_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_1_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_2_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_2_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_3_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_3_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_4_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_4_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_5_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_5_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_6_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_6_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_7_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_7_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_8_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_8_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_9_s_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_9_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_10_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_10_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_10_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_11_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_11_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_11_1_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_12_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_12_U.t_read | ~AESL_inst_example.edge_index_cpy2_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_example.edge_index_cpy2_V_12_1_U.t_read | ((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_2[2] = dl_detect_out ? proc_dep_vld_vec_2_reg[2] : (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_2[3] = dl_detect_out ? proc_dep_vld_vec_2_reg[3] : (((AESL_inst_example.clone_vector_1_U0_ap_ready_count[0]) & AESL_inst_example.clone_vector_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[11 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[23 : 12] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign in_chan_dep_vld_vec_2[2] = dep_chan_vld_3_2;
    assign in_chan_dep_data_vec_2[35 : 24] = dep_chan_data_3_2;
    assign token_in_vec_2[2] = token_3_2;
    assign in_chan_dep_vld_vec_2[3] = dep_chan_vld_5_2;
    assign in_chan_dep_data_vec_2[47 : 36] = dep_chan_data_5_2;
    assign token_in_vec_2[3] = token_5_2;
    assign dep_chan_vld_2_3 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_3 = out_chan_dep_data_2;
    assign token_2_3 = token_out_vec_2[0];
    assign dep_chan_vld_2_5 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_5 = out_chan_dep_data_2;
    assign token_2_5 = token_out_vec_2[1];
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[2];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[2];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[3];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[3];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$clone_vector_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$clone_vector_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$clone_vector_U0$ap_idle <= AESL_inst_example.clone_vector_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.clone_vector_U0
    AESL_deadlock_detect_unit #(12, 3, 3, 3) AESL_deadlock_detect_unit_3 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (~AESL_inst_example.edge_index_cpy1_0_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_0_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_0_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_0_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_1_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_1_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_1_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_1_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_2_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_2_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_2_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_2_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_3_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_3_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_3_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_3_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_4_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_4_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_4_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_4_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_5_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_5_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_5_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_5_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_6_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_6_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_6_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_6_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_7_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_7_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_7_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_7_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_8_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_8_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_8_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_8_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_9_0_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_9_0_U.i_write | ~AESL_inst_example.edge_index_cpy1_9_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_9_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_10_s_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_10_s_U.i_write | ~AESL_inst_example.edge_index_cpy1_10_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_10_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_11_s_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_11_s_U.i_write | ~AESL_inst_example.edge_index_cpy1_11_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_11_1_U.i_write | ~AESL_inst_example.edge_index_cpy1_12_s_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_12_s_U.i_write | ~AESL_inst_example.edge_index_cpy1_12_1_U.t_empty_n & (AESL_inst_example.clone_vector_U0.ap_ready | AESL_inst_example.clone_vector_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy1_12_1_U.i_write);
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (~AESL_inst_example.edge_index_cpy3_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_0_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_0_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_0_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_1_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_1_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_1_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_2_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_2_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_2_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_3_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_3_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_3_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_4_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_4_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_4_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_5_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_5_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_5_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_6_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_6_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_6_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_7_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_7_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_7_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_8_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_8_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_8_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_9_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_9_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_9_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_10_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_10_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_10_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_11_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_11_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_11_3_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_12_1_U.t_read | ~AESL_inst_example.edge_index_cpy3_V_12_3_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy3_V_12_3_U.t_read);
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (~AESL_inst_example.edge_index_cpy4_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_0_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_0_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_1_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_1_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_2_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_2_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_3_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_3_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_4_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_4_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_5_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_5_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_6_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_6_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_7_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_7_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_8_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_8_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_9_s_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_9_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_10_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_10_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_10_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_11_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_11_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_11_1_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_12_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_12_U.t_read | ~AESL_inst_example.edge_index_cpy4_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_example.edge_index_cpy4_V_12_1_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_2_3;
    assign in_chan_dep_data_vec_3[11 : 0] = dep_chan_data_2_3;
    assign token_in_vec_3[0] = token_2_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_7_3;
    assign in_chan_dep_data_vec_3[23 : 12] = dep_chan_data_7_3;
    assign token_in_vec_3[1] = token_7_3;
    assign in_chan_dep_vld_vec_3[2] = dep_chan_vld_11_3;
    assign in_chan_dep_data_vec_3[35 : 24] = dep_chan_data_11_3;
    assign token_in_vec_3[2] = token_11_3;
    assign dep_chan_vld_3_2 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_2 = out_chan_dep_data_3;
    assign token_3_2 = token_out_vec_3[0];
    assign dep_chan_vld_3_7 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_7 = out_chan_dep_data_3;
    assign token_3_7 = token_out_vec_3[1];
    assign dep_chan_vld_3_11 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_11 = out_chan_dep_data_3;
    assign token_3_11 = token_out_vec_3[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Loop_edge_choose_ver_1_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Loop_edge_choose_ver_1_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Loop_edge_choose_ver_1_U0$ap_idle <= AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Loop_edge_choose_ver_1_U0
    AESL_deadlock_detect_unit #(12, 4, 2, 2) AESL_deadlock_detect_unit_4 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (~AESL_inst_example.node_attr_cpy1_V_0_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_0_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_1_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_1_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_2_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_2_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_3_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_3_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_4_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_4_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_5_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_5_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_6_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_6_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_7_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_7_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_8_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_8_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_9_0_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_9_0_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_10_s_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_10_s_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_0_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_1_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_2_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_3_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_4_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_5_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_6_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_7_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_8_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_9_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_10_1_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_0_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_1_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_2_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_3_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_4_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_5_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_6_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_7_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_8_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_9_2_U.i_write | ~AESL_inst_example.node_attr_cpy1_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy1_V_10_2_U.i_write);
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_0_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_12_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_12_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_2_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_2_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_3_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_3_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_4_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_4_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_5_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_5_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_6_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_6_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_7_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_7_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_8_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_8_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_9_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_9_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_15_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_15_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_18_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_18_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_21_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_21_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_0_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_0_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_12_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_12_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_2_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_2_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_3_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_3_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_4_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_4_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_5_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_5_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_6_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_6_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_7_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_7_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_8_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_8_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_9_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_9_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_15_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_15_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_18_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_18_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_21_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_21_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_0_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_0_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_13_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_13_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_2_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_2_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_3_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_3_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_4_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_4_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_5_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_5_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_6_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_6_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_7_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_7_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_8_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_8_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_9_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_9_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_16_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_16_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_19_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_19_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_22_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_22_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_0_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_0_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_13_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_13_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_2_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_2_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_3_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_3_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_4_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_4_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_5_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_5_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_6_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_6_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_7_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_7_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_8_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_8_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_9_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_9_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_16_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_16_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_19_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_19_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_22_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_22_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_0_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_0_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_14_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_14_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_2_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_2_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_3_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_3_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_4_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_4_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_5_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_5_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_6_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_6_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_7_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_7_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_8_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_8_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_9_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_9_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_17_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_17_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_20_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_20_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_23_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_s_mat_1_23_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_0_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_0_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_14_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_14_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_2_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_2_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_3_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_3_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_4_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_4_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_5_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_5_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_6_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_6_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_7_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_7_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_8_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_8_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_9_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_9_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_17_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_17_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_20_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_20_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_23_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_1_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_example.node_attr_1D_r_mat_1_23_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_1_4;
    assign in_chan_dep_data_vec_4[11 : 0] = dep_chan_data_1_4;
    assign token_in_vec_4[0] = token_1_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_5_4;
    assign in_chan_dep_data_vec_4[23 : 12] = dep_chan_data_5_4;
    assign token_in_vec_4[1] = token_5_4;
    assign dep_chan_vld_4_1 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_1 = out_chan_dep_data_4;
    assign token_4_1 = token_out_vec_4[0];
    assign dep_chan_vld_4_5 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_5 = out_chan_dep_data_4;
    assign token_4_5 = token_out_vec_4[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Loop_edge_compute_lo_1_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Loop_edge_compute_lo_1_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Loop_edge_compute_lo_1_U0$ap_idle <= AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Loop_edge_compute_lo_1_U0
    AESL_deadlock_detect_unit #(12, 5, 5, 5) AESL_deadlock_detect_unit_5 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (~AESL_inst_example.edge_index_cpy2_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_0_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_0_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_1_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_1_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_2_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_2_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_3_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_3_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_4_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_4_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_5_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_5_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_6_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_6_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_7_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_7_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_8_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_8_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_9_s_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_9_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_10_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_10_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_11_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_11_1_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_12_U.i_write | ~AESL_inst_example.edge_index_cpy2_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy2_V_12_1_U.i_write | ((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_1_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (~AESL_inst_example.node_attr_1D_s_mat_0_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_0_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_0_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_0_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_0_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_0_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_12_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_12_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_13_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_13_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_13_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_13_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_14_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_14_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_14_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_14_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_2_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_2_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_2_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_2_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_2_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_2_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_3_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_3_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_3_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_3_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_3_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_3_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_4_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_4_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_4_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_4_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_4_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_4_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_5_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_5_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_5_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_5_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_5_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_5_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_6_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_6_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_6_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_6_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_6_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_6_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_7_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_7_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_7_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_7_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_7_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_7_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_8_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_8_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_8_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_8_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_8_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_8_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_9_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_9_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_9_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_9_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_9_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_9_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_15_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_15_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_15_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_15_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_16_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_16_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_16_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_16_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_17_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_17_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_17_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_17_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_18_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_18_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_18_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_18_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_19_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_19_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_19_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_19_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_20_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_20_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_20_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_20_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_21_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_21_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_21_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_21_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_22_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_22_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_22_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_22_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_23_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_23_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_23_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_23_U.i_write);
    assign proc_dep_vld_vec_5[2] = dl_detect_out ? proc_dep_vld_vec_5_reg[2] : (~AESL_inst_example.layer7_out_0_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_0_V_U.t_read | ~AESL_inst_example.layer7_out_0_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_1_V_U.t_read | ~AESL_inst_example.layer7_out_0_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_2_V_U.t_read | ~AESL_inst_example.layer7_out_0_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_0_3_V_U.t_read | ~AESL_inst_example.layer7_out_1_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_0_V_U.t_read | ~AESL_inst_example.layer7_out_1_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_1_V_U.t_read | ~AESL_inst_example.layer7_out_1_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_2_V_U.t_read | ~AESL_inst_example.layer7_out_1_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_1_3_V_U.t_read | ~AESL_inst_example.layer7_out_2_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_0_V_U.t_read | ~AESL_inst_example.layer7_out_2_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_1_V_U.t_read | ~AESL_inst_example.layer7_out_2_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_2_V_U.t_read | ~AESL_inst_example.layer7_out_2_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_2_3_V_U.t_read | ~AESL_inst_example.layer7_out_3_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_0_V_U.t_read | ~AESL_inst_example.layer7_out_3_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_1_V_U.t_read | ~AESL_inst_example.layer7_out_3_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_2_V_U.t_read | ~AESL_inst_example.layer7_out_3_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_3_3_V_U.t_read | ~AESL_inst_example.layer7_out_4_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_0_V_U.t_read | ~AESL_inst_example.layer7_out_4_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_1_V_U.t_read | ~AESL_inst_example.layer7_out_4_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_2_V_U.t_read | ~AESL_inst_example.layer7_out_4_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_4_3_V_U.t_read | ~AESL_inst_example.layer7_out_5_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_0_V_U.t_read | ~AESL_inst_example.layer7_out_5_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_1_V_U.t_read | ~AESL_inst_example.layer7_out_5_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_2_V_U.t_read | ~AESL_inst_example.layer7_out_5_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_5_3_V_U.t_read | ~AESL_inst_example.layer7_out_6_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_0_V_U.t_read | ~AESL_inst_example.layer7_out_6_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_1_V_U.t_read | ~AESL_inst_example.layer7_out_6_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_2_V_U.t_read | ~AESL_inst_example.layer7_out_6_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_6_3_V_U.t_read | ~AESL_inst_example.layer7_out_7_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_0_V_U.t_read | ~AESL_inst_example.layer7_out_7_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_1_V_U.t_read | ~AESL_inst_example.layer7_out_7_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_2_V_U.t_read | ~AESL_inst_example.layer7_out_7_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_7_3_V_U.t_read | ~AESL_inst_example.layer7_out_8_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_0_V_U.t_read | ~AESL_inst_example.layer7_out_8_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_1_V_U.t_read | ~AESL_inst_example.layer7_out_8_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_2_V_U.t_read | ~AESL_inst_example.layer7_out_8_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_8_3_V_U.t_read | ~AESL_inst_example.layer7_out_9_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_0_V_U.t_read | ~AESL_inst_example.layer7_out_9_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_1_V_U.t_read | ~AESL_inst_example.layer7_out_9_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_2_V_U.t_read | ~AESL_inst_example.layer7_out_9_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_9_3_V_U.t_read | ~AESL_inst_example.layer7_out_10_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_0_V_U.t_read | ~AESL_inst_example.layer7_out_10_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_1_V_U.t_read | ~AESL_inst_example.layer7_out_10_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_2_V_U.t_read | ~AESL_inst_example.layer7_out_10_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_10_3_V_U.t_read | ~AESL_inst_example.layer7_out_11_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_0_V_U.t_read | ~AESL_inst_example.layer7_out_11_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_1_V_U.t_read | ~AESL_inst_example.layer7_out_11_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_2_V_U.t_read | ~AESL_inst_example.layer7_out_11_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_11_3_V_U.t_read | ~AESL_inst_example.layer7_out_12_0_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_0_V_U.t_read | ~AESL_inst_example.layer7_out_12_1_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_1_V_U.t_read | ~AESL_inst_example.layer7_out_12_2_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_2_V_U.t_read | ~AESL_inst_example.layer7_out_12_3_V_U.i_full_n & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_example.layer7_out_12_3_V_U.t_read);
    assign proc_dep_vld_vec_5[3] = dl_detect_out ? proc_dep_vld_vec_5_reg[3] : (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.Block_proc_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_5[4] = dl_detect_out ? proc_dep_vld_vec_5_reg[4] : (((AESL_inst_example.Loop_edge_compute_lo_1_U0_ap_ready_count[0]) & AESL_inst_example.Loop_edge_compute_lo_1_U0.ap_idle & ~(AESL_inst_example.clone_vector_3_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_0_5;
    assign in_chan_dep_data_vec_5[11 : 0] = dep_chan_data_0_5;
    assign token_in_vec_5[0] = token_0_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_1_5;
    assign in_chan_dep_data_vec_5[23 : 12] = dep_chan_data_1_5;
    assign token_in_vec_5[1] = token_1_5;
    assign in_chan_dep_vld_vec_5[2] = dep_chan_vld_2_5;
    assign in_chan_dep_data_vec_5[35 : 24] = dep_chan_data_2_5;
    assign token_in_vec_5[2] = token_2_5;
    assign in_chan_dep_vld_vec_5[3] = dep_chan_vld_4_5;
    assign in_chan_dep_data_vec_5[47 : 36] = dep_chan_data_4_5;
    assign token_in_vec_5[3] = token_4_5;
    assign in_chan_dep_vld_vec_5[4] = dep_chan_vld_6_5;
    assign in_chan_dep_data_vec_5[59 : 48] = dep_chan_data_6_5;
    assign token_in_vec_5[4] = token_6_5;
    assign dep_chan_vld_5_2 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_2 = out_chan_dep_data_5;
    assign token_5_2 = token_out_vec_5[0];
    assign dep_chan_vld_5_4 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_4 = out_chan_dep_data_5;
    assign token_5_4 = token_out_vec_5[1];
    assign dep_chan_vld_5_6 = out_chan_dep_vld_vec_5[2];
    assign dep_chan_data_5_6 = out_chan_dep_data_5;
    assign token_5_6 = token_out_vec_5[2];
    assign dep_chan_vld_5_0 = out_chan_dep_vld_vec_5[3];
    assign dep_chan_data_5_0 = out_chan_dep_data_5;
    assign token_5_0 = token_out_vec_5[3];
    assign dep_chan_vld_5_1 = out_chan_dep_vld_vec_5[4];
    assign dep_chan_data_5_1 = out_chan_dep_data_5;
    assign token_5_1 = token_out_vec_5[4];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$clone_vector_2_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$clone_vector_2_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$clone_vector_2_U0$ap_idle <= AESL_inst_example.clone_vector_2_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.clone_vector_2_U0
    AESL_deadlock_detect_unit #(12, 6, 3, 3) AESL_deadlock_detect_unit_6 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (~AESL_inst_example.layer7_out_0_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_0_V_U.i_write | ~AESL_inst_example.layer7_out_0_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_1_V_U.i_write | ~AESL_inst_example.layer7_out_0_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_2_V_U.i_write | ~AESL_inst_example.layer7_out_0_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_0_3_V_U.i_write | ~AESL_inst_example.layer7_out_1_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_0_V_U.i_write | ~AESL_inst_example.layer7_out_1_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_1_V_U.i_write | ~AESL_inst_example.layer7_out_1_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_2_V_U.i_write | ~AESL_inst_example.layer7_out_1_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_1_3_V_U.i_write | ~AESL_inst_example.layer7_out_2_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_0_V_U.i_write | ~AESL_inst_example.layer7_out_2_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_1_V_U.i_write | ~AESL_inst_example.layer7_out_2_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_2_V_U.i_write | ~AESL_inst_example.layer7_out_2_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_2_3_V_U.i_write | ~AESL_inst_example.layer7_out_3_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_0_V_U.i_write | ~AESL_inst_example.layer7_out_3_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_1_V_U.i_write | ~AESL_inst_example.layer7_out_3_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_2_V_U.i_write | ~AESL_inst_example.layer7_out_3_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_3_3_V_U.i_write | ~AESL_inst_example.layer7_out_4_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_0_V_U.i_write | ~AESL_inst_example.layer7_out_4_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_1_V_U.i_write | ~AESL_inst_example.layer7_out_4_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_2_V_U.i_write | ~AESL_inst_example.layer7_out_4_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_4_3_V_U.i_write | ~AESL_inst_example.layer7_out_5_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_0_V_U.i_write | ~AESL_inst_example.layer7_out_5_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_1_V_U.i_write | ~AESL_inst_example.layer7_out_5_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_2_V_U.i_write | ~AESL_inst_example.layer7_out_5_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_5_3_V_U.i_write | ~AESL_inst_example.layer7_out_6_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_0_V_U.i_write | ~AESL_inst_example.layer7_out_6_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_1_V_U.i_write | ~AESL_inst_example.layer7_out_6_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_2_V_U.i_write | ~AESL_inst_example.layer7_out_6_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_6_3_V_U.i_write | ~AESL_inst_example.layer7_out_7_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_0_V_U.i_write | ~AESL_inst_example.layer7_out_7_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_1_V_U.i_write | ~AESL_inst_example.layer7_out_7_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_2_V_U.i_write | ~AESL_inst_example.layer7_out_7_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_7_3_V_U.i_write | ~AESL_inst_example.layer7_out_8_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_0_V_U.i_write | ~AESL_inst_example.layer7_out_8_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_1_V_U.i_write | ~AESL_inst_example.layer7_out_8_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_2_V_U.i_write | ~AESL_inst_example.layer7_out_8_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_8_3_V_U.i_write | ~AESL_inst_example.layer7_out_9_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_0_V_U.i_write | ~AESL_inst_example.layer7_out_9_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_1_V_U.i_write | ~AESL_inst_example.layer7_out_9_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_2_V_U.i_write | ~AESL_inst_example.layer7_out_9_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_9_3_V_U.i_write | ~AESL_inst_example.layer7_out_10_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_0_V_U.i_write | ~AESL_inst_example.layer7_out_10_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_1_V_U.i_write | ~AESL_inst_example.layer7_out_10_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_2_V_U.i_write | ~AESL_inst_example.layer7_out_10_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_10_3_V_U.i_write | ~AESL_inst_example.layer7_out_11_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_0_V_U.i_write | ~AESL_inst_example.layer7_out_11_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_1_V_U.i_write | ~AESL_inst_example.layer7_out_11_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_2_V_U.i_write | ~AESL_inst_example.layer7_out_11_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_11_3_V_U.i_write | ~AESL_inst_example.layer7_out_12_0_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_0_V_U.i_write | ~AESL_inst_example.layer7_out_12_1_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_1_V_U.i_write | ~AESL_inst_example.layer7_out_12_2_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_2_V_U.i_write | ~AESL_inst_example.layer7_out_12_3_V_U.t_empty_n & (AESL_inst_example.clone_vector_2_U0.ap_ready | AESL_inst_example.clone_vector_2_U0.ap_idle) & ~AESL_inst_example.layer7_out_12_3_V_U.i_write);
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (~AESL_inst_example.layer7_out_cpy1_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_0_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_0_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_0_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_0_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_0_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_0_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_1_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_1_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_2_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_2_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_3_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_3_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_4_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_4_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_5_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_5_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_6_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_6_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_7_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_7_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_8_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_8_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_s_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_9_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_9_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_10_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_10_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_11_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_11_7_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_1_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_2_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_3_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_4_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_4_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_5_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_5_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_6_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_6_U.t_read | ~AESL_inst_example.layer7_out_cpy1_V_12_7_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy1_V_12_7_U.t_read);
    assign proc_dep_vld_vec_6[2] = dl_detect_out ? proc_dep_vld_vec_6_reg[2] : (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_0_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_0_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_0_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_0_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_1_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_1_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_1_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_1_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_1_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_2_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_2_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_2_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_2_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_2_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_3_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_3_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_3_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_3_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_3_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_4_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_4_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_4_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_4_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_4_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_5_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_5_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_5_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_5_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_5_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_6_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_6_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_6_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_6_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_6_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_7_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_7_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_7_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_7_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_7_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_8_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_8_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_8_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_8_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_8_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_9_s_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_s_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_9_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_9_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_9_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_9_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_10_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_10_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_10_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_10_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_10_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_11_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_11_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_11_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_11_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_11_3_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_12_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_12_1_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_1_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_12_2_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_2_U.t_read | ~AESL_inst_example.layer7_out_cpy2_V_12_3_U.i_full_n & AESL_inst_example.clone_vector_2_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_example.layer7_out_cpy2_V_12_3_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_5_6;
    assign in_chan_dep_data_vec_6[11 : 0] = dep_chan_data_5_6;
    assign token_in_vec_6[0] = token_5_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_7_6;
    assign in_chan_dep_data_vec_6[23 : 12] = dep_chan_data_7_6;
    assign token_in_vec_6[1] = token_7_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_11_6;
    assign in_chan_dep_data_vec_6[35 : 24] = dep_chan_data_11_6;
    assign token_in_vec_6[2] = token_11_6;
    assign dep_chan_vld_6_5 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_5 = out_chan_dep_data_6;
    assign token_6_5 = token_out_vec_6[0];
    assign dep_chan_vld_6_7 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_7 = out_chan_dep_data_6;
    assign token_6_7 = token_out_vec_6[1];
    assign dep_chan_vld_6_11 = out_chan_dep_vld_vec_6[2];
    assign dep_chan_data_6_11 = out_chan_dep_data_6;
    assign token_6_11 = token_out_vec_6[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Loop_fetch_loop_proc_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Loop_fetch_loop_proc_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Loop_fetch_loop_proc_U0$ap_idle <= AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Loop_fetch_loop_proc_U0
    AESL_deadlock_detect_unit #(12, 7, 3, 3) AESL_deadlock_detect_unit_7 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (~AESL_inst_example.edge_attr_aggr_0_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_0_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_0_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_1_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_1_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_2_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_2_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_3_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_3_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_4_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_4_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_5_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_5_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_6_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_6_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_7_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_7_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_8_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_8_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_9_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_9_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_10_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_10_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_11_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_11_3_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_0_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_0_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_0_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_0_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_0_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_1_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_1_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_1_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_1_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_2_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_2_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_2_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_2_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_3_1_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_1_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_3_2_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_2_U.t_read | ~AESL_inst_example.edge_attr_aggr_12_3_3_U.i_full_n & AESL_inst_example.Loop_fetch_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_example.edge_attr_aggr_12_3_3_U.t_read);
    assign proc_dep_vld_vec_7[1] = dl_detect_out ? proc_dep_vld_vec_7_reg[1] : (~AESL_inst_example.edge_index_cpy3_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_0_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_0_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_0_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_1_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_1_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_1_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_2_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_2_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_2_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_3_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_3_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_3_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_4_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_4_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_4_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_5_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_5_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_5_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_6_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_6_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_6_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_7_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_7_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_7_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_8_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_8_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_8_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_9_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_9_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_9_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_10_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_10_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_10_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_11_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_11_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_11_3_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_12_1_U.i_write | ~AESL_inst_example.edge_index_cpy3_V_12_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy3_V_12_3_U.i_write);
    assign proc_dep_vld_vec_7[2] = dl_detect_out ? proc_dep_vld_vec_7_reg[2] : (~AESL_inst_example.layer7_out_cpy1_V_12_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_12_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_12_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_12_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_4_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_4_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_5_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_5_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_6_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_6_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_7_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_7_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_12_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_12_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_12_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_12_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_11_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_11_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_10_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_10_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_9_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_9_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_8_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_8_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_7_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_7_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_6_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_6_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_5_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_5_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_4_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_4_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_3_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_3_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_2_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_2_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_1_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_1_3_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_s_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_1_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_2_U.i_write | ~AESL_inst_example.layer7_out_cpy1_V_0_3_U.t_empty_n & (AESL_inst_example.Loop_fetch_loop_proc_U0.ap_ready | AESL_inst_example.Loop_fetch_loop_proc_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy1_V_0_3_U.i_write);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_3_7;
    assign in_chan_dep_data_vec_7[11 : 0] = dep_chan_data_3_7;
    assign token_in_vec_7[0] = token_3_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_6_7;
    assign in_chan_dep_data_vec_7[23 : 12] = dep_chan_data_6_7;
    assign token_in_vec_7[1] = token_6_7;
    assign in_chan_dep_vld_vec_7[2] = dep_chan_vld_8_7;
    assign in_chan_dep_data_vec_7[35 : 24] = dep_chan_data_8_7;
    assign token_in_vec_7[2] = token_8_7;
    assign dep_chan_vld_7_8 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_8 = out_chan_dep_data_7;
    assign token_7_8 = token_out_vec_7[0];
    assign dep_chan_vld_7_3 = out_chan_dep_vld_vec_7[1];
    assign dep_chan_data_7_3 = out_chan_dep_data_7;
    assign token_7_3 = token_out_vec_7[1];
    assign dep_chan_vld_7_6 = out_chan_dep_vld_vec_7[2];
    assign dep_chan_data_7_6 = out_chan_dep_data_7;
    assign token_7_6 = token_out_vec_7[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Loop_out_loop_proc_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Loop_out_loop_proc_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Loop_out_loop_proc_U0$ap_idle <= AESL_inst_example.Loop_out_loop_proc_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Loop_out_loop_proc_U0
    AESL_deadlock_detect_unit #(12, 8, 2, 2) AESL_deadlock_detect_unit_8 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (~AESL_inst_example.edge_attr_aggr_0_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_0_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_0_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_1_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_2_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_3_1_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_1_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_0_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_1_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_2_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_3_2_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_2_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_0_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_0_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_1_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_1_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_2_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_2_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_3_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_3_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_4_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_4_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_5_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_5_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_6_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_6_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_7_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_7_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_8_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_8_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_9_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_9_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_10_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_10_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_11_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_11_3_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_0_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_0_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_1_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_1_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_2_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_2_3_U.i_write | ~AESL_inst_example.edge_attr_aggr_12_3_3_U.t_empty_n & (AESL_inst_example.Loop_out_loop_proc_U0.ap_ready | AESL_inst_example.Loop_out_loop_proc_U0.ap_idle) & ~AESL_inst_example.edge_attr_aggr_12_3_3_U.i_write);
    assign proc_dep_vld_vec_8[1] = dl_detect_out ? proc_dep_vld_vec_8_reg[1] : (~AESL_inst_example.layer9_out_1_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_0_V_U.t_read | ~AESL_inst_example.layer9_out_2_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_0_V_U.t_read | ~AESL_inst_example.layer9_out_3_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_0_V_U.t_read | ~AESL_inst_example.layer9_out_4_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_0_V_U.t_read | ~AESL_inst_example.layer9_out_5_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_0_V_U.t_read | ~AESL_inst_example.layer9_out_6_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_0_V_U.t_read | ~AESL_inst_example.layer9_out_7_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_0_V_U.t_read | ~AESL_inst_example.layer9_out_8_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_0_V_U.t_read | ~AESL_inst_example.layer9_out_9_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_0_V_U.t_read | ~AESL_inst_example.layer9_out_10_0_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_0_V_U.t_read | ~AESL_inst_example.layer9_out_1_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_1_V_U.t_read | ~AESL_inst_example.layer9_out_2_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_1_V_U.t_read | ~AESL_inst_example.layer9_out_3_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_1_V_U.t_read | ~AESL_inst_example.layer9_out_4_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_1_V_U.t_read | ~AESL_inst_example.layer9_out_5_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_1_V_U.t_read | ~AESL_inst_example.layer9_out_6_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_1_V_U.t_read | ~AESL_inst_example.layer9_out_7_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_1_V_U.t_read | ~AESL_inst_example.layer9_out_8_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_1_V_U.t_read | ~AESL_inst_example.layer9_out_9_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_1_V_U.t_read | ~AESL_inst_example.layer9_out_10_1_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_1_V_U.t_read | ~AESL_inst_example.layer9_out_1_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_2_V_U.t_read | ~AESL_inst_example.layer9_out_2_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_2_V_U.t_read | ~AESL_inst_example.layer9_out_3_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_2_V_U.t_read | ~AESL_inst_example.layer9_out_4_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_2_V_U.t_read | ~AESL_inst_example.layer9_out_5_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_2_V_U.t_read | ~AESL_inst_example.layer9_out_6_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_2_V_U.t_read | ~AESL_inst_example.layer9_out_7_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_2_V_U.t_read | ~AESL_inst_example.layer9_out_8_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_2_V_U.t_read | ~AESL_inst_example.layer9_out_9_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_2_V_U.t_read | ~AESL_inst_example.layer9_out_10_2_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_2_V_U.t_read | ~AESL_inst_example.layer9_out_1_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_1_3_V_U.t_read | ~AESL_inst_example.layer9_out_2_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_2_3_V_U.t_read | ~AESL_inst_example.layer9_out_3_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_3_3_V_U.t_read | ~AESL_inst_example.layer9_out_4_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_4_3_V_U.t_read | ~AESL_inst_example.layer9_out_5_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_5_3_V_U.t_read | ~AESL_inst_example.layer9_out_6_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_6_3_V_U.t_read | ~AESL_inst_example.layer9_out_7_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_7_3_V_U.t_read | ~AESL_inst_example.layer9_out_8_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_8_3_V_U.t_read | ~AESL_inst_example.layer9_out_9_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_9_3_V_U.t_read | ~AESL_inst_example.layer9_out_10_3_V_U.i_full_n & AESL_inst_example.Loop_out_loop_proc_U0.ap_done & deadlock_detector.ap_done_reg_7 & ~AESL_inst_example.layer9_out_10_3_V_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_7_8;
    assign in_chan_dep_data_vec_8[11 : 0] = dep_chan_data_7_8;
    assign token_in_vec_8[0] = token_7_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_9_8;
    assign in_chan_dep_data_vec_8[23 : 12] = dep_chan_data_9_8;
    assign token_in_vec_8[1] = token_9_8;
    assign dep_chan_vld_8_7 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_7 = out_chan_dep_data_8;
    assign token_8_7 = token_out_vec_8[0];
    assign dep_chan_vld_8_9 = out_chan_dep_vld_vec_8[1];
    assign dep_chan_data_8_9 = out_chan_dep_data_8;
    assign token_8_9 = token_out_vec_8[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Loop_node_compute_lo_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Loop_node_compute_lo_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Loop_node_compute_lo_U0$ap_idle <= AESL_inst_example.Loop_node_compute_lo_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Loop_node_compute_lo_U0
    AESL_deadlock_detect_unit #(12, 9, 3, 3) AESL_deadlock_detect_unit_9 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (~AESL_inst_example.node_attr_cpy2_V_0_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_0_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_0_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_0_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_1_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_1_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_1_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_1_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_2_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_2_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_2_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_2_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_3_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_3_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_3_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_3_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_4_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_4_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_4_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_4_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_5_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_5_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_5_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_5_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_6_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_6_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_6_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_6_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_7_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_7_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_7_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_7_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_8_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_8_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_8_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_8_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_9_0_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_9_0_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_9_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_9_2_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_10_s_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_10_s_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_10_1_U.i_write | ~AESL_inst_example.node_attr_cpy2_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_cpy2_V_10_2_U.i_write);
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (~AESL_inst_example.layer10_out_0_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_0_0_V_U.t_read | ~AESL_inst_example.layer10_out_0_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_0_1_V_U.t_read | ~AESL_inst_example.layer10_out_0_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_0_2_V_U.t_read | ~AESL_inst_example.layer10_out_1_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_1_0_V_U.t_read | ~AESL_inst_example.layer10_out_1_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_1_1_V_U.t_read | ~AESL_inst_example.layer10_out_1_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_1_2_V_U.t_read | ~AESL_inst_example.layer10_out_2_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_2_0_V_U.t_read | ~AESL_inst_example.layer10_out_2_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_2_1_V_U.t_read | ~AESL_inst_example.layer10_out_2_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_2_2_V_U.t_read | ~AESL_inst_example.layer10_out_3_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_3_0_V_U.t_read | ~AESL_inst_example.layer10_out_3_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_3_1_V_U.t_read | ~AESL_inst_example.layer10_out_3_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_3_2_V_U.t_read | ~AESL_inst_example.layer10_out_4_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_4_0_V_U.t_read | ~AESL_inst_example.layer10_out_4_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_4_1_V_U.t_read | ~AESL_inst_example.layer10_out_4_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_4_2_V_U.t_read | ~AESL_inst_example.layer10_out_5_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_5_0_V_U.t_read | ~AESL_inst_example.layer10_out_5_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_5_1_V_U.t_read | ~AESL_inst_example.layer10_out_5_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_5_2_V_U.t_read | ~AESL_inst_example.layer10_out_6_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_6_0_V_U.t_read | ~AESL_inst_example.layer10_out_6_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_6_1_V_U.t_read | ~AESL_inst_example.layer10_out_6_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_6_2_V_U.t_read | ~AESL_inst_example.layer10_out_7_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_7_0_V_U.t_read | ~AESL_inst_example.layer10_out_7_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_7_1_V_U.t_read | ~AESL_inst_example.layer10_out_7_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_7_2_V_U.t_read | ~AESL_inst_example.layer10_out_8_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_8_0_V_U.t_read | ~AESL_inst_example.layer10_out_8_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_8_1_V_U.t_read | ~AESL_inst_example.layer10_out_8_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_8_2_V_U.t_read | ~AESL_inst_example.layer10_out_9_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_9_0_V_U.t_read | ~AESL_inst_example.layer10_out_9_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_9_1_V_U.t_read | ~AESL_inst_example.layer10_out_9_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_9_2_V_U.t_read | ~AESL_inst_example.layer10_out_10_0_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_10_0_V_U.t_read | ~AESL_inst_example.layer10_out_10_1_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_10_1_V_U.t_read | ~AESL_inst_example.layer10_out_10_2_V_U.i_full_n & AESL_inst_example.Loop_node_compute_lo_U0.ap_done & deadlock_detector.ap_done_reg_8 & ~AESL_inst_example.layer10_out_10_2_V_U.t_read);
    assign proc_dep_vld_vec_9[2] = dl_detect_out ? proc_dep_vld_vec_9_reg[2] : (~AESL_inst_example.layer9_out_1_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_0_V_U.i_write | ~AESL_inst_example.layer9_out_1_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_1_V_U.i_write | ~AESL_inst_example.layer9_out_1_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_2_V_U.i_write | ~AESL_inst_example.layer9_out_1_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_1_3_V_U.i_write | ~AESL_inst_example.layer9_out_2_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_0_V_U.i_write | ~AESL_inst_example.layer9_out_2_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_1_V_U.i_write | ~AESL_inst_example.layer9_out_2_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_2_V_U.i_write | ~AESL_inst_example.layer9_out_2_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_2_3_V_U.i_write | ~AESL_inst_example.layer9_out_3_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_0_V_U.i_write | ~AESL_inst_example.layer9_out_3_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_1_V_U.i_write | ~AESL_inst_example.layer9_out_3_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_2_V_U.i_write | ~AESL_inst_example.layer9_out_3_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_3_3_V_U.i_write | ~AESL_inst_example.layer9_out_4_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_0_V_U.i_write | ~AESL_inst_example.layer9_out_4_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_1_V_U.i_write | ~AESL_inst_example.layer9_out_4_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_2_V_U.i_write | ~AESL_inst_example.layer9_out_4_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_4_3_V_U.i_write | ~AESL_inst_example.layer9_out_5_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_0_V_U.i_write | ~AESL_inst_example.layer9_out_5_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_1_V_U.i_write | ~AESL_inst_example.layer9_out_5_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_2_V_U.i_write | ~AESL_inst_example.layer9_out_5_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_5_3_V_U.i_write | ~AESL_inst_example.layer9_out_6_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_0_V_U.i_write | ~AESL_inst_example.layer9_out_6_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_1_V_U.i_write | ~AESL_inst_example.layer9_out_6_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_2_V_U.i_write | ~AESL_inst_example.layer9_out_6_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_6_3_V_U.i_write | ~AESL_inst_example.layer9_out_7_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_0_V_U.i_write | ~AESL_inst_example.layer9_out_7_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_1_V_U.i_write | ~AESL_inst_example.layer9_out_7_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_2_V_U.i_write | ~AESL_inst_example.layer9_out_7_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_7_3_V_U.i_write | ~AESL_inst_example.layer9_out_8_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_0_V_U.i_write | ~AESL_inst_example.layer9_out_8_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_1_V_U.i_write | ~AESL_inst_example.layer9_out_8_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_2_V_U.i_write | ~AESL_inst_example.layer9_out_8_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_8_3_V_U.i_write | ~AESL_inst_example.layer9_out_9_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_0_V_U.i_write | ~AESL_inst_example.layer9_out_9_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_1_V_U.i_write | ~AESL_inst_example.layer9_out_9_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_2_V_U.i_write | ~AESL_inst_example.layer9_out_9_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_9_3_V_U.i_write | ~AESL_inst_example.layer9_out_10_0_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_0_V_U.i_write | ~AESL_inst_example.layer9_out_10_1_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_1_V_U.i_write | ~AESL_inst_example.layer9_out_10_2_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_2_V_U.i_write | ~AESL_inst_example.layer9_out_10_3_V_U.t_empty_n & (AESL_inst_example.Loop_node_compute_lo_U0.ap_ready | AESL_inst_example.Loop_node_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer9_out_10_3_V_U.i_write);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_1_9;
    assign in_chan_dep_data_vec_9[11 : 0] = dep_chan_data_1_9;
    assign token_in_vec_9[0] = token_1_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_8_9;
    assign in_chan_dep_data_vec_9[23 : 12] = dep_chan_data_8_9;
    assign token_in_vec_9[1] = token_8_9;
    assign in_chan_dep_vld_vec_9[2] = dep_chan_vld_10_9;
    assign in_chan_dep_data_vec_9[35 : 24] = dep_chan_data_10_9;
    assign token_in_vec_9[2] = token_10_9;
    assign dep_chan_vld_9_1 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_1 = out_chan_dep_data_9;
    assign token_9_1 = token_out_vec_9[0];
    assign dep_chan_vld_9_10 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_10 = out_chan_dep_data_9;
    assign token_9_10 = token_out_vec_9[1];
    assign dep_chan_vld_9_8 = out_chan_dep_vld_vec_9[2];
    assign dep_chan_data_9_8 = out_chan_dep_data_9;
    assign token_9_8 = token_out_vec_9[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Loop_edge_choose_ver_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Loop_edge_choose_ver_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Loop_edge_choose_ver_U0$ap_idle <= AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Loop_edge_choose_ver_U0
    AESL_deadlock_detect_unit #(12, 10, 2, 2) AESL_deadlock_detect_unit_10 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (~AESL_inst_example.layer10_out_0_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_0_0_V_U.i_write | ~AESL_inst_example.layer10_out_1_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_1_0_V_U.i_write | ~AESL_inst_example.layer10_out_2_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_2_0_V_U.i_write | ~AESL_inst_example.layer10_out_3_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_3_0_V_U.i_write | ~AESL_inst_example.layer10_out_4_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_4_0_V_U.i_write | ~AESL_inst_example.layer10_out_5_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_5_0_V_U.i_write | ~AESL_inst_example.layer10_out_6_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_6_0_V_U.i_write | ~AESL_inst_example.layer10_out_7_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_7_0_V_U.i_write | ~AESL_inst_example.layer10_out_8_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_8_0_V_U.i_write | ~AESL_inst_example.layer10_out_9_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_9_0_V_U.i_write | ~AESL_inst_example.layer10_out_10_0_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_10_0_V_U.i_write | ~AESL_inst_example.layer10_out_0_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_0_1_V_U.i_write | ~AESL_inst_example.layer10_out_1_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_1_1_V_U.i_write | ~AESL_inst_example.layer10_out_2_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_2_1_V_U.i_write | ~AESL_inst_example.layer10_out_3_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_3_1_V_U.i_write | ~AESL_inst_example.layer10_out_4_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_4_1_V_U.i_write | ~AESL_inst_example.layer10_out_5_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_5_1_V_U.i_write | ~AESL_inst_example.layer10_out_6_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_6_1_V_U.i_write | ~AESL_inst_example.layer10_out_7_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_7_1_V_U.i_write | ~AESL_inst_example.layer10_out_8_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_8_1_V_U.i_write | ~AESL_inst_example.layer10_out_9_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_9_1_V_U.i_write | ~AESL_inst_example.layer10_out_10_1_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_10_1_V_U.i_write | ~AESL_inst_example.layer10_out_0_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_0_2_V_U.i_write | ~AESL_inst_example.layer10_out_1_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_1_2_V_U.i_write | ~AESL_inst_example.layer10_out_2_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_2_2_V_U.i_write | ~AESL_inst_example.layer10_out_3_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_3_2_V_U.i_write | ~AESL_inst_example.layer10_out_4_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_4_2_V_U.i_write | ~AESL_inst_example.layer10_out_5_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_5_2_V_U.i_write | ~AESL_inst_example.layer10_out_6_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_6_2_V_U.i_write | ~AESL_inst_example.layer10_out_7_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_7_2_V_U.i_write | ~AESL_inst_example.layer10_out_8_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_8_2_V_U.i_write | ~AESL_inst_example.layer10_out_9_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_9_2_V_U.i_write | ~AESL_inst_example.layer10_out_10_2_V_U.t_empty_n & (AESL_inst_example.Loop_edge_choose_ver_U0.ap_ready | AESL_inst_example.Loop_edge_choose_ver_U0.ap_idle) & ~AESL_inst_example.layer10_out_10_2_V_U.i_write);
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (~AESL_inst_example.node_attr_1D_s_mat_0_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_0_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_6_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_7_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_8_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_9_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_3_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_6_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_9_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_0_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_0_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_6_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_7_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_8_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_9_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_3_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_3_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_6_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_6_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_9_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_9_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_0_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_0_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_2_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_2_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_3_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_3_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_4_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_4_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_5_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_5_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_6_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_6_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_7_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_7_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_8_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_8_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_9_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_9_1_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_4_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_7_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_10_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_10_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_0_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_0_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_2_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_2_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_3_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_3_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_4_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_4_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_5_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_5_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_6_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_6_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_7_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_7_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_8_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_8_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_9_1_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_9_1_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_4_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_4_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_7_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_7_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_10_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_10_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_0_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_0_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_2_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_2_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_3_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_3_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_4_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_4_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_5_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_5_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_6_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_6_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_7_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_7_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_8_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_8_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_9_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_9_2_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_5_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_8_U.t_read | ~AESL_inst_example.node_attr_1D_s_mat_1_11_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_s_mat_1_11_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_0_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_0_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_2_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_2_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_3_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_3_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_4_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_4_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_5_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_5_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_6_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_6_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_7_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_7_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_8_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_8_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_9_2_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_9_2_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_5_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_5_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_8_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_8_U.t_read | ~AESL_inst_example.node_attr_1D_r_mat_1_11_U.i_full_n & AESL_inst_example.Loop_edge_choose_ver_U0.ap_done & deadlock_detector.ap_done_reg_9 & ~AESL_inst_example.node_attr_1D_r_mat_1_11_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_9_10;
    assign in_chan_dep_data_vec_10[11 : 0] = dep_chan_data_9_10;
    assign token_in_vec_10[0] = token_9_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_11_10;
    assign in_chan_dep_data_vec_10[23 : 12] = dep_chan_data_11_10;
    assign token_in_vec_10[1] = token_11_10;
    assign dep_chan_vld_10_9 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_9 = out_chan_dep_data_10;
    assign token_10_9 = token_out_vec_10[0];
    assign dep_chan_vld_10_11 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_11 = out_chan_dep_data_10;
    assign token_10_11 = token_out_vec_10[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_example$Loop_edge_compute_lo_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_example$Loop_edge_compute_lo_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_example$Loop_edge_compute_lo_U0$ap_idle <= AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle;
        end
    end
    // Process: AESL_inst_example.Loop_edge_compute_lo_U0
    AESL_deadlock_detect_unit #(12, 11, 3, 3) AESL_deadlock_detect_unit_11 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_11),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_11),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_11),
        .token_in_vec(token_in_vec_11),
        .dl_detect_in(dl_detect_out),
        .origin(origin[11]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_11),
        .out_chan_dep_data(out_chan_dep_data_11),
        .token_out_vec(token_out_vec_11),
        .dl_detect_out(dl_in_vec[11]));

    assign proc_dep_vld_vec_11[0] = dl_detect_out ? proc_dep_vld_vec_11_reg[0] : (~AESL_inst_example.layer7_out_cpy2_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_0_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_0_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_1_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_1_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_2_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_2_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_3_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_3_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_4_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_4_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_5_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_5_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_6_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_6_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_7_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_7_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_8_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_8_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_s_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_9_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_9_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_10_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_10_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_10_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_11_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_11_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_11_3_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_1_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_12_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_2_U.i_write | ~AESL_inst_example.layer7_out_cpy2_V_12_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.layer7_out_cpy2_V_12_3_U.i_write);
    assign proc_dep_vld_vec_11[1] = dl_detect_out ? proc_dep_vld_vec_11_reg[1] : (~AESL_inst_example.edge_index_cpy4_V_0_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_0_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_0_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_1_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_1_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_1_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_2_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_2_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_2_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_3_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_3_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_3_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_4_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_4_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_4_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_5_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_5_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_5_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_6_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_6_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_6_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_7_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_7_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_7_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_8_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_8_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_8_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_9_s_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_9_s_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_9_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_10_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_10_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_10_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_11_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_11_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_11_1_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_12_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_12_U.i_write | ~AESL_inst_example.edge_index_cpy4_V_12_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.edge_index_cpy4_V_12_1_U.i_write);
    assign proc_dep_vld_vec_11[2] = dl_detect_out ? proc_dep_vld_vec_11_reg[2] : (~AESL_inst_example.node_attr_1D_s_mat_0_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_0_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_0_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_0_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_0_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_0_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_2_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_2_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_2_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_2_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_3_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_3_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_3_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_3_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_4_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_4_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_4_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_4_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_5_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_5_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_5_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_5_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_6_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_6_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_6_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_6_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_7_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_7_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_7_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_7_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_8_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_8_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_8_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_8_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_1_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_9_1_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_1_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_9_2_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_9_2_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_9_2_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_3_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_3_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_3_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_4_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_4_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_4_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_5_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_5_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_5_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_6_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_6_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_6_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_7_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_7_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_7_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_8_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_8_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_8_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_9_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_9_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_9_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_10_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_10_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_10_U.i_write | ~AESL_inst_example.node_attr_1D_s_mat_1_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_s_mat_1_11_U.i_write | ~AESL_inst_example.node_attr_1D_r_mat_1_11_U.t_empty_n & (AESL_inst_example.Loop_edge_compute_lo_U0.ap_ready | AESL_inst_example.Loop_edge_compute_lo_U0.ap_idle) & ~AESL_inst_example.node_attr_1D_r_mat_1_11_U.i_write);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_11_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_11_reg <= proc_dep_vld_vec_11;
        end
    end
    assign in_chan_dep_vld_vec_11[0] = dep_chan_vld_3_11;
    assign in_chan_dep_data_vec_11[11 : 0] = dep_chan_data_3_11;
    assign token_in_vec_11[0] = token_3_11;
    assign in_chan_dep_vld_vec_11[1] = dep_chan_vld_6_11;
    assign in_chan_dep_data_vec_11[23 : 12] = dep_chan_data_6_11;
    assign token_in_vec_11[1] = token_6_11;
    assign in_chan_dep_vld_vec_11[2] = dep_chan_vld_10_11;
    assign in_chan_dep_data_vec_11[35 : 24] = dep_chan_data_10_11;
    assign token_in_vec_11[2] = token_10_11;
    assign dep_chan_vld_11_6 = out_chan_dep_vld_vec_11[0];
    assign dep_chan_data_11_6 = out_chan_dep_data_11;
    assign token_11_6 = token_out_vec_11[0];
    assign dep_chan_vld_11_3 = out_chan_dep_vld_vec_11[1];
    assign dep_chan_data_11_3 = out_chan_dep_data_11;
    assign token_11_3 = token_out_vec_11[1];
    assign dep_chan_vld_11_10 = out_chan_dep_vld_vec_11[2];
    assign dep_chan_data_11_10 = out_chan_dep_data_11;
    assign token_11_10 = token_out_vec_11[2];


    AESL_deadlock_report_unit #(12) AESL_deadlock_report_unit_inst (
        .reset(reset),
        .clock(clock),
        .dl_in_vec(dl_in_vec),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
